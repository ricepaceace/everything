
module Decision ( ap_clk, ap_rst_n, s_axi_AXILiteS_AWVALID, 
        s_axi_AXILiteS_AWREADY, s_axi_AXILiteS_AWADDR, s_axi_AXILiteS_WVALID, 
        s_axi_AXILiteS_WREADY, s_axi_AXILiteS_WDATA, s_axi_AXILiteS_WSTRB, 
        s_axi_AXILiteS_ARVALID, s_axi_AXILiteS_ARREADY, s_axi_AXILiteS_ARADDR, 
        s_axi_AXILiteS_RVALID, s_axi_AXILiteS_RREADY, s_axi_AXILiteS_RDATA, 
        s_axi_AXILiteS_RRESP, s_axi_AXILiteS_BVALID, s_axi_AXILiteS_BREADY, 
        s_axi_AXILiteS_BRESP, interrupt );
  input [6:0] s_axi_AXILiteS_AWADDR;
  input [31:0] s_axi_AXILiteS_WDATA;
  input [3:0] s_axi_AXILiteS_WSTRB;
  input [6:0] s_axi_AXILiteS_ARADDR;
  output [31:0] s_axi_AXILiteS_RDATA;
  output [1:0] s_axi_AXILiteS_RRESP;
  output [1:0] s_axi_AXILiteS_BRESP;
  input ap_clk, ap_rst_n, s_axi_AXILiteS_AWVALID, s_axi_AXILiteS_WVALID,
         s_axi_AXILiteS_ARVALID, s_axi_AXILiteS_RREADY, s_axi_AXILiteS_BREADY;
  output s_axi_AXILiteS_AWREADY, s_axi_AXILiteS_WREADY, s_axi_AXILiteS_ARREADY,
         s_axi_AXILiteS_RVALID, s_axi_AXILiteS_BVALID, interrupt;
  wire   \tmp_s_reg_1578[0] , \recentVBools_data_q0[0] ,
         \recentVBools_data_q1[0] , \tmp_12_reg_1694[0] ,
         \recentABools_data_q0[0] , \recentABools_data_q1[0] , ap_start,
         \reset_A_V[0] , \reset_V_V[0] , \reset_params_V[0] , N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         \last_sample_is_A_V[0] , \last_sample_is_V_V[0] ,
         \last_sample_is_V_V_loc_2_reg_358[0] , \tmp_13_reg_1725[0] ,
         \tmp_8_reg_1630[0] , \tmp_19_reg_409[0] , \not_tmp_i_i2_reg_1745[0] ,
         \not_tmp_i_i4_reg_1650[0] , \tmp_i3_reg_1674[0] ,
         \recentABools_data_load_reg_1700[0] , \tmp_22_reg_1772[0] ,
         \tmp_25_reg_1777[0] , \recentVBools_data_load_reg_1584[0] ,
         \toReturn_5_reg_1655[0] , \toReturn_6_reg_1660[0] ,
         \toReturn_7_reg_1750[0] , \toReturn_8_reg_1755[0] , N461, N466, N472,
         i_fu_607_p2_31, p_1_cast_fu_1031_p1_31, p_cast_fu_688_p1_31, N495,
         N496, N497, N498, N499, N500, N502, N503, N505, N512, N513,
         toReturn_1_fu_1395_p3_12, \toReturn_1_fu_1395_p3[7] ,
         \dp_cluster_0/N985 , \dp_cluster_0/N984 , \dp_cluster_0/N983 ,
         \dp_cluster_0/N982 , \dp_cluster_0/N981 , \dp_cluster_0/N980 ,
         \dp_cluster_0/N979 , \dp_cluster_0/N978 , \dp_cluster_0/N977 ,
         \dp_cluster_0/N976 , \dp_cluster_0/N975 , \dp_cluster_0/N974 ,
         \dp_cluster_0/N973 , \dp_cluster_0/N972 , \dp_cluster_0/N971 ,
         \dp_cluster_0/N970 , \dp_cluster_0/N969 , \dp_cluster_0/N968 ,
         \dp_cluster_0/N967 , \dp_cluster_0/N966 , \dp_cluster_0/N965 ,
         \dp_cluster_0/N964 , \dp_cluster_0/N963 , \dp_cluster_0/N962 ,
         \dp_cluster_0/N961 , \dp_cluster_0/N960 , \dp_cluster_0/N959 ,
         \dp_cluster_0/N958 , \dp_cluster_0/N957 , \dp_cluster_0/N956 ,
         \dp_cluster_0/N955 , \dp_cluster_0/N954 , \dp_cluster_1/N953 ,
         \dp_cluster_1/N952 , \dp_cluster_1/N951 , \dp_cluster_1/N950 ,
         \dp_cluster_1/N949 , \dp_cluster_1/N948 , \dp_cluster_1/N947 ,
         \dp_cluster_1/N946 , \dp_cluster_1/N945 , \dp_cluster_1/N944 ,
         \dp_cluster_1/N943 , \dp_cluster_1/N942 , \dp_cluster_1/N941 ,
         \dp_cluster_1/N940 , \dp_cluster_1/N939 , \dp_cluster_1/N938 ,
         \dp_cluster_1/N937 , \dp_cluster_1/N936 , \dp_cluster_1/N935 ,
         \dp_cluster_1/N934 , \dp_cluster_1/N933 , \dp_cluster_1/N932 ,
         \dp_cluster_1/N931 , \dp_cluster_1/N930 , \dp_cluster_1/N929 ,
         \dp_cluster_1/N928 , \dp_cluster_1/N927 , \dp_cluster_1/N926 ,
         \dp_cluster_1/N925 , \dp_cluster_1/N924 , \dp_cluster_1/N923 ,
         \dp_cluster_1/N922 ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[0] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[10] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[11] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[12] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[13] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[14] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[15] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[16] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[17] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[18] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[19] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[1] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[20] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[21] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[22] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[23] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[24] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[25] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[26] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[27] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[28] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[29] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[2] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[30] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[31] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[3] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[4] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[5] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[6] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[7] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[8] ,
         \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[9] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[0] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[10] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[11] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[12] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[13] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[14] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[15] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[16] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[17] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[18] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[19] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[1] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[20] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[21] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[22] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[23] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[24] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[25] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[26] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[27] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[28] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[29] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[2] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[30] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[31] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[3] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[4] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[5] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[6] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[7] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[8] ,
         \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[9] , n264,
         n265, n266, n267, n268, n269, n272, n276, n277, n278, n282, n285,
         n286, n287, n288, n289, n290, n298, n299, n302, n305, n306, n307,
         n308, n309, n310, n311, n312, n318, n319, n322, n325, n326, n327,
         n328, n329, n330, n338, n339, n342, n345, n346, n347, n349, n350,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n367, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n397, n398, n399,
         n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410,
         n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
         n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432,
         n433, n436, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n478, n483, n486, n489, n491,
         n493, n494, n496, n497, n499, n500, n502, n503, n505, n506, n508,
         n509, n511, n512, n514, n515, n517, n518, n520, n521, n523, n524,
         n526, n527, n529, n530, n532, n533, n535, n536, n538, n539, n541,
         n542, n544, n545, n547, n548, n550, n551, n553, n554, n556, n557,
         n559, n560, n562, n563, n565, n566, n568, n569, n571, n572, n574,
         n575, n577, n578, n580, n581, n583, n584, n585, n588, n590, n591,
         n593, n594, n596, n597, n599, n600, n602, n603, n605, n606, n608,
         n609, n611, n612, n614, n615, n617, n618, n620, n621, n623, n624,
         n626, n627, n629, n630, n632, n633, n635, n636, n638, n639, n641,
         n642, n644, n645, n647, n648, n650, n651, n653, n654, n656, n657,
         n659, n660, n662, n663, n665, n666, n668, n669, n671, n672, n674,
         n675, n677, n678, n680, n681, n683, n684, n685, n686, n688, n689,
         n691, n692, n694, n696, n698, n700, n702, n703, n705, n706, n708,
         n710, n712, n714, n716, n717, n719, n720, n722, n723, n725, n727,
         n729, n730, n732, n733, n735, n737, n739, n741, n743, n744, n746,
         n747, n749, n751, n753, n755, n757, n758, n760, n761, n763, n764,
         n766, n767, n769, n770, n772, n773, n775, n777, n779, n781, n783,
         n784, n786, n788, n790, n792, n793, n794, n795, n798, n799, n800,
         n803, n806, n807, n808, n809, n813, n816, n817, n818, n821, n824,
         n825, n826, n827, n830, n833, n834, n836, n837, n838, n839, n840,
         n841, n842, n843, n850, n851, n854, n857, n858, n859, n860, n861,
         n862, n869, n870, n873, n877, n880, n882, n884, n885, n886, n888,
         n890, n891, n892, n894, n896, n897, n899, n901, n902, n903, n904,
         n905, n907, n909, n911, n913, n914, n915, n916, n918, n920, n921,
         n922, n924, n925, n926, n927, n928, n930, n932, n933, n934, n936,
         n938, n940, n942, n943, n944, n945, n946, n947, n948, n949, n951,
         n953, n954, n955, n957, n959, n961, n962, n963, n964, n965, n966,
         n967, n968, n970, n972, n973, n975, n976, n978, n979, n981, n983,
         n985, n987, n989, n990, n992, n993, n995, n997, n999, n1001, n1003,
         n1004, n1006, n1007, n1009, n1011, n1013, n1014, n1016, n1017, n1019,
         n1021, n1023, n1025, n1027, n1028, n1030, n1031, n1033, n1034, n1036,
         n1037, n1039, n1041, n1043, n1045, n1047, n1048, n1050, n1051, n1053,
         n1054, n1056, n1057, n1059, n1060, n1062, n1064, n1066, n1068, n1069,
         n1071, n1073, n1075, n1076, n1078, n1080, n1082, n1084, n1086, n1088,
         n1090, n1092, n1094, n1096, n1098, n1100, n1102, n1104, n1106, n1108,
         n1110, n1112, n1114, n1116, n1118, n1120, n1122, n1124, n1126, n1128,
         n1130, n1132, n1134, n1136, n1138, n1140, n1142, n1144, n1146, n1148,
         n1150, n1152, n1154, n1156, n1158, n1160, n1162, n1164, n1166, n1168,
         n1170, n1172, n1174, n1176, n1178, n1180, n1182, n1184, n1186, n1188,
         n1190, n1192, n1194, n1196, n1198, n1200, n1202, n1204, n1206, n1208,
         n1210, n1212, n1213, n1216, n1218, n1219, n1221, n1223, n1224, n1226,
         n1228, n1229, n1230, n1231, n1232, n1234, n1235, n1236, n1237, n1238,
         n1245, n1246, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1263, n1264, n1267, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1281, n1282, n1284, n1285, n1286, n1287, n1288,
         n1289, n1291, n1292, n1294, n1295, n1297, n1298, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1319, n1320, n1322, n1323, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1334, n1336, n1338,
         n1340, n1342, n1344, n1346, n1348, n1350, n1352, n1354, n1356, n1358,
         n1360, n1362, n1364, n1366, n1368, n1370, n1372, n1374, n1376, n1378,
         n1380, n1382, n1384, n1386, n1388, n1390, n1392, n1394, n1396, n1398,
         n1400, n1401, n1404, n1406, n1408, n1410, n1412, n1414, n1416, n1418,
         n1420, n1422, n1424, n1426, n1428, n1430, n1432, n1434, n1436, n1438,
         n1440, n1442, n1444, n1446, n1448, n1450, n1452, n1454, n1456, n1458,
         n1460, n1462, n1464, n1466, n1468, n1469, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1485, n1486, n1489, n1492, n1493, n1494,
         n1495, n1496, n1497, n1504, n1505, n1508, n1512, n1513, n1514, n1515,
         n1516, n1517, n1520, n1521, n1522, n1525, n1528, n1529, n1530, n1531,
         n1535, n1538, n1539, n1540, n1543, n1546, n1547, n1548, n1549, n1552,
         n1556, n1558, n1560, n1561, n1562, n1564, n1566, n1567, n1568, n1570,
         n1572, n1573, n1575, n1577, n1578, n1579, n1580, n1581, n1583, n1585,
         n1587, n1589, n1590, n1591, n1592, n1594, n1596, n1597, n1598, n1600,
         n1601, n1602, n1603, n1604, n1606, n1608, n1609, n1610, n1612, n1614,
         n1616, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1627,
         n1629, n1630, n1631, n1633, n1635, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1646, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1664, n1665, n1668, n1672, n1673, n1674,
         n1675, n1676, n1677, n1685, n1686, n1689, n1693, n1695, n1696, n1699,
         n1701, n1702, n1703, n1704, n1706, n1708, n1709, n1711, n1712, n1714,
         n1715, n1717, n1718, n1720, n1721, n1723, n1724, n1726, n1727, n1729,
         n1730, n1732, n1733, n1735, n1736, n1738, n1739, n1741, n1742, n1744,
         n1745, n1747, n1748, n1750, n1751, n1753, n1754, n1756, n1757, n1759,
         n1760, n1762, n1763, n1765, n1766, n1768, n1769, n1771, n1772, n1774,
         n1775, n1777, n1778, n1780, n1781, n1783, n1784, n1786, n1787, n1789,
         n1790, n1792, n1794, n1796, n1798, n1800, n1801, n1802, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1831, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1843, n1845, n1847, n1848, n1849, n1851, n1853,
         n1854, n1855, n1856, n1857, n1859, n1861, n1863, n1865, n1867, n1869,
         n1872, n1874, n1876, n1878, n1880, n1882, n1884, n1886, n1888, n1890,
         n1892, n1894, n1896, n1898, n1900, n1902, n1904, n1906, n1908, n1910,
         n1912, n1914, n1916, n1918, n1920, n1922, n1924, n1926, n1928, n1930,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1980, n1983, n1986,
         n1988, n2017, n2018, n2020, n2022, n2024, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2190, n2192, n2193, n2194, n2195, n2196,
         n2198, n2199, n2200, n2201, n2202, n2203, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2237, n2238, n2239, n2240,
         n2241, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2294, n2296, n2298, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2336,
         n2340, n2342, n2344, n2346, n2348, n2350, n2352, n2354, n2356, n2358,
         n2360, n2362, n2364, n2366, n2368, n2370, n2372, n2374, n2376, n2378,
         n2380, n2382, n2384, n2386, n2388, n2390, n2392, n2394, n2396, n2398,
         n2400, n2401, n2402, n2403, n2406, n2408, n2410, n2412, n2414, n2416,
         n2418, n2420, n2422, n2424, n2426, n2428, n2430, n2432, n2434, n2436,
         n2438, n2440, n2442, n2444, n2446, n2448, n2450, n2452, n2454, n2456,
         n2458, n2460, n2462, n2464, n2466, n2468, n2470, n2472, n2474, n2476,
         n2478, n2480, n2482, n2484, n2486, n2488, n2490, n2492, n2494, n2496,
         n2498, n2500, n2502, n2504, n2506, n2508, n2510, n2512, n2514, n2516,
         n2518, n2520, n2522, n2524, n2526, n2528, n2530, n2532, n2533, n2534,
         n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543, n2544,
         n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553, n2554,
         n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563, n2564,
         n2565, n2566, n2567, n2571, n2574, n2576, n2578, n2580, n2582, n2584,
         n2586, n2588, n2590, n2592, n2594, n2596, n2598, n2600, n2602, n2604,
         n2606, n2608, n2610, n2612, n2614, n2616, n2618, n2620, n2622, n2624,
         n2626, n2628, n2630, n2632, n2634, n2636, n2638, n2640, n2642, n2644,
         n2646, n2648, n2650, n2652, n2654, n2656, n2658, n2660, n2662, n2664,
         n2666, n2668, n2670, n2672, n2674, n2676, n2678, n2680, n2682, n2684,
         n2686, n2688, n2690, n2692, n2694, n2696, n2698, n2699, n2700, n2701,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2787, n2789, n2791, n2793, n2794, n2795, n2797,
         n2801, n2803, n2805, n2807, n2809, n2811, n2813, n2815, n2817, n2819,
         n2821, n2823, n2825, n2827, n2829, n2831, n2833, n2835, n2837, n2839,
         n2841, n2843, n2845, n2847, n2849, n2851, n2853, n2855, n2857, n2859,
         n2861, n2862, n2863, n2864, n2865, n2867, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2936, n2938, n2940, n2942, n2944, n2946, n2948, n2950,
         n2952, n2954, n2956, n2958, n2960, n2962, n2964, n2966, n2968, n2970,
         n2972, n2974, n2976, n2978, n2980, n2982, n2984, n2986, n2988, n2990,
         n2992, n2994, n2996, n2998, n2999, n3000, n3001, n3002, n3003, n3004,
         n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014,
         n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024,
         n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034,
         n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044,
         n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054,
         n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3064, n3066,
         n3068, n3070, n3072, n3074, n3076, n3078, n3080, n3082, n3084, n3086,
         n3088, n3090, n3092, n3094, n3096, n3098, n3100, n3102, n3104, n3106,
         n3108, n3110, n3112, n3114, n3116, n3118, n3120, n3122, n3124, n3126,
         n3127, n3128, n3130, n3132, n3133, n3134, n3136, n3138, n3139, n3140,
         n3142, n3144, n3145, n3146, n3149, n3151, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616,
         n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626,
         n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636,
         n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646,
         n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656,
         n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666,
         n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676,
         n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686,
         n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696,
         n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706,
         n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716,
         n3717, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4214,
         n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224,
         n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234,
         n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244,
         n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254,
         n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264,
         n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274,
         n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304,
         n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314,
         n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324,
         n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334,
         n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344,
         n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354,
         n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364,
         n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374,
         n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384,
         n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394,
         n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404,
         n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414,
         n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424,
         n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434,
         n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444,
         n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454,
         n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464,
         n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474,
         n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484,
         n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494,
         n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504,
         n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514,
         n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524,
         n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554,
         n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564,
         n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574,
         n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584,
         n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594,
         n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634,
         n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644,
         n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674,
         n4675, n4676, n4677, n4678, n4679, n4680,
         \Decision_AXILiteS_s_axi_U/n873 , \Decision_AXILiteS_s_axi_U/n871 ,
         \Decision_AXILiteS_s_axi_U/n870 , \Decision_AXILiteS_s_axi_U/n869 ,
         \Decision_AXILiteS_s_axi_U/n868 , \Decision_AXILiteS_s_axi_U/n867 ,
         \Decision_AXILiteS_s_axi_U/n866 , \Decision_AXILiteS_s_axi_U/n865 ,
         \Decision_AXILiteS_s_axi_U/n863 , \Decision_AXILiteS_s_axi_U/n862 ,
         \Decision_AXILiteS_s_axi_U/n861 , \Decision_AXILiteS_s_axi_U/n860 ,
         \Decision_AXILiteS_s_axi_U/n859 , \Decision_AXILiteS_s_axi_U/n858 ,
         \Decision_AXILiteS_s_axi_U/n857 , \Decision_AXILiteS_s_axi_U/n856 ,
         \Decision_AXILiteS_s_axi_U/n855 , \Decision_AXILiteS_s_axi_U/n854 ,
         \Decision_AXILiteS_s_axi_U/n853 , \Decision_AXILiteS_s_axi_U/n852 ,
         \Decision_AXILiteS_s_axi_U/n851 , \Decision_AXILiteS_s_axi_U/n850 ,
         \Decision_AXILiteS_s_axi_U/n849 , \Decision_AXILiteS_s_axi_U/n848 ,
         \Decision_AXILiteS_s_axi_U/n847 , \Decision_AXILiteS_s_axi_U/n846 ,
         \Decision_AXILiteS_s_axi_U/n845 , \Decision_AXILiteS_s_axi_U/n844 ,
         \Decision_AXILiteS_s_axi_U/n843 , \Decision_AXILiteS_s_axi_U/n842 ,
         \Decision_AXILiteS_s_axi_U/n841 , \Decision_AXILiteS_s_axi_U/n840 ,
         \Decision_AXILiteS_s_axi_U/n839 , \Decision_AXILiteS_s_axi_U/n838 ,
         \Decision_AXILiteS_s_axi_U/n837 , \Decision_AXILiteS_s_axi_U/n836 ,
         \Decision_AXILiteS_s_axi_U/n835 , \Decision_AXILiteS_s_axi_U/n834 ,
         \Decision_AXILiteS_s_axi_U/n833 , \Decision_AXILiteS_s_axi_U/n832 ,
         \Decision_AXILiteS_s_axi_U/n831 , \Decision_AXILiteS_s_axi_U/n830 ,
         \Decision_AXILiteS_s_axi_U/n829 , \Decision_AXILiteS_s_axi_U/n828 ,
         \Decision_AXILiteS_s_axi_U/n827 , \Decision_AXILiteS_s_axi_U/n826 ,
         \Decision_AXILiteS_s_axi_U/n825 , \Decision_AXILiteS_s_axi_U/n824 ,
         \Decision_AXILiteS_s_axi_U/n823 , \Decision_AXILiteS_s_axi_U/n822 ,
         \Decision_AXILiteS_s_axi_U/n821 , \Decision_AXILiteS_s_axi_U/n820 ,
         \Decision_AXILiteS_s_axi_U/n819 , \Decision_AXILiteS_s_axi_U/n818 ,
         \Decision_AXILiteS_s_axi_U/n817 , \Decision_AXILiteS_s_axi_U/n816 ,
         \Decision_AXILiteS_s_axi_U/n815 , \Decision_AXILiteS_s_axi_U/n814 ,
         \Decision_AXILiteS_s_axi_U/n813 , \Decision_AXILiteS_s_axi_U/n812 ,
         \Decision_AXILiteS_s_axi_U/n811 , \Decision_AXILiteS_s_axi_U/n810 ,
         \Decision_AXILiteS_s_axi_U/n809 , \Decision_AXILiteS_s_axi_U/n808 ,
         \Decision_AXILiteS_s_axi_U/n807 , \Decision_AXILiteS_s_axi_U/n806 ,
         \Decision_AXILiteS_s_axi_U/n805 , \Decision_AXILiteS_s_axi_U/n804 ,
         \Decision_AXILiteS_s_axi_U/n803 , \Decision_AXILiteS_s_axi_U/n802 ,
         \Decision_AXILiteS_s_axi_U/n801 , \Decision_AXILiteS_s_axi_U/n800 ,
         \Decision_AXILiteS_s_axi_U/n799 , \Decision_AXILiteS_s_axi_U/n798 ,
         \Decision_AXILiteS_s_axi_U/n797 , \Decision_AXILiteS_s_axi_U/n796 ,
         \Decision_AXILiteS_s_axi_U/n795 , \Decision_AXILiteS_s_axi_U/n794 ,
         \Decision_AXILiteS_s_axi_U/n793 , \Decision_AXILiteS_s_axi_U/n792 ,
         \Decision_AXILiteS_s_axi_U/n791 , \Decision_AXILiteS_s_axi_U/n790 ,
         \Decision_AXILiteS_s_axi_U/n789 , \Decision_AXILiteS_s_axi_U/n788 ,
         \Decision_AXILiteS_s_axi_U/n787 , \Decision_AXILiteS_s_axi_U/n786 ,
         \Decision_AXILiteS_s_axi_U/n785 , \Decision_AXILiteS_s_axi_U/n784 ,
         \Decision_AXILiteS_s_axi_U/n783 , \Decision_AXILiteS_s_axi_U/n782 ,
         \Decision_AXILiteS_s_axi_U/n781 , \Decision_AXILiteS_s_axi_U/n780 ,
         \Decision_AXILiteS_s_axi_U/n779 , \Decision_AXILiteS_s_axi_U/n778 ,
         \Decision_AXILiteS_s_axi_U/n777 , \Decision_AXILiteS_s_axi_U/n776 ,
         \Decision_AXILiteS_s_axi_U/n775 , \Decision_AXILiteS_s_axi_U/n774 ,
         \Decision_AXILiteS_s_axi_U/n773 , \Decision_AXILiteS_s_axi_U/n772 ,
         \Decision_AXILiteS_s_axi_U/n771 , \Decision_AXILiteS_s_axi_U/n770 ,
         \Decision_AXILiteS_s_axi_U/n769 , \Decision_AXILiteS_s_axi_U/n768 ,
         \Decision_AXILiteS_s_axi_U/n767 , \Decision_AXILiteS_s_axi_U/n766 ,
         \Decision_AXILiteS_s_axi_U/n765 , \Decision_AXILiteS_s_axi_U/n764 ,
         \Decision_AXILiteS_s_axi_U/n763 , \Decision_AXILiteS_s_axi_U/n762 ,
         \Decision_AXILiteS_s_axi_U/n761 , \Decision_AXILiteS_s_axi_U/n760 ,
         \Decision_AXILiteS_s_axi_U/n759 , \Decision_AXILiteS_s_axi_U/n758 ,
         \Decision_AXILiteS_s_axi_U/n757 , \Decision_AXILiteS_s_axi_U/n756 ,
         \Decision_AXILiteS_s_axi_U/n755 , \Decision_AXILiteS_s_axi_U/n754 ,
         \Decision_AXILiteS_s_axi_U/n753 , \Decision_AXILiteS_s_axi_U/n752 ,
         \Decision_AXILiteS_s_axi_U/n751 , \Decision_AXILiteS_s_axi_U/n750 ,
         \Decision_AXILiteS_s_axi_U/n749 , \Decision_AXILiteS_s_axi_U/n748 ,
         \Decision_AXILiteS_s_axi_U/n747 , \Decision_AXILiteS_s_axi_U/n746 ,
         \Decision_AXILiteS_s_axi_U/n745 , \Decision_AXILiteS_s_axi_U/n744 ,
         \Decision_AXILiteS_s_axi_U/n743 , \Decision_AXILiteS_s_axi_U/n742 ,
         \Decision_AXILiteS_s_axi_U/n741 , \Decision_AXILiteS_s_axi_U/n740 ,
         \Decision_AXILiteS_s_axi_U/n739 , \Decision_AXILiteS_s_axi_U/n738 ,
         \Decision_AXILiteS_s_axi_U/n737 , \Decision_AXILiteS_s_axi_U/n736 ,
         \Decision_AXILiteS_s_axi_U/n735 , \Decision_AXILiteS_s_axi_U/n734 ,
         \Decision_AXILiteS_s_axi_U/n733 , \Decision_AXILiteS_s_axi_U/n732 ,
         \Decision_AXILiteS_s_axi_U/n731 , \Decision_AXILiteS_s_axi_U/n730 ,
         \Decision_AXILiteS_s_axi_U/n729 , \Decision_AXILiteS_s_axi_U/n728 ,
         \Decision_AXILiteS_s_axi_U/n727 , \Decision_AXILiteS_s_axi_U/n726 ,
         \Decision_AXILiteS_s_axi_U/n725 , \Decision_AXILiteS_s_axi_U/n724 ,
         \Decision_AXILiteS_s_axi_U/n723 , \Decision_AXILiteS_s_axi_U/n722 ,
         \Decision_AXILiteS_s_axi_U/n721 , \Decision_AXILiteS_s_axi_U/n720 ,
         \Decision_AXILiteS_s_axi_U/n719 , \Decision_AXILiteS_s_axi_U/n718 ,
         \Decision_AXILiteS_s_axi_U/n717 , \Decision_AXILiteS_s_axi_U/n716 ,
         \Decision_AXILiteS_s_axi_U/n715 , \Decision_AXILiteS_s_axi_U/n714 ,
         \Decision_AXILiteS_s_axi_U/n713 , \Decision_AXILiteS_s_axi_U/n712 ,
         \Decision_AXILiteS_s_axi_U/n711 , \Decision_AXILiteS_s_axi_U/n710 ,
         \Decision_AXILiteS_s_axi_U/n709 , \Decision_AXILiteS_s_axi_U/n708 ,
         \Decision_AXILiteS_s_axi_U/n707 , \Decision_AXILiteS_s_axi_U/n706 ,
         \Decision_AXILiteS_s_axi_U/n705 , \Decision_AXILiteS_s_axi_U/n704 ,
         \Decision_AXILiteS_s_axi_U/n703 , \Decision_AXILiteS_s_axi_U/n702 ,
         \Decision_AXILiteS_s_axi_U/n701 , \Decision_AXILiteS_s_axi_U/n700 ,
         \Decision_AXILiteS_s_axi_U/n699 , \Decision_AXILiteS_s_axi_U/n698 ,
         \Decision_AXILiteS_s_axi_U/n697 , \Decision_AXILiteS_s_axi_U/n696 ,
         \Decision_AXILiteS_s_axi_U/n695 , \Decision_AXILiteS_s_axi_U/n694 ,
         \Decision_AXILiteS_s_axi_U/n693 , \Decision_AXILiteS_s_axi_U/n692 ,
         \Decision_AXILiteS_s_axi_U/n691 , \Decision_AXILiteS_s_axi_U/n690 ,
         \Decision_AXILiteS_s_axi_U/n689 , \Decision_AXILiteS_s_axi_U/n688 ,
         \Decision_AXILiteS_s_axi_U/n687 , \Decision_AXILiteS_s_axi_U/n686 ,
         \Decision_AXILiteS_s_axi_U/n685 , \Decision_AXILiteS_s_axi_U/n684 ,
         \Decision_AXILiteS_s_axi_U/n683 , \Decision_AXILiteS_s_axi_U/n682 ,
         \Decision_AXILiteS_s_axi_U/n681 , \Decision_AXILiteS_s_axi_U/n680 ,
         \Decision_AXILiteS_s_axi_U/n679 , \Decision_AXILiteS_s_axi_U/n678 ,
         \Decision_AXILiteS_s_axi_U/n677 , \Decision_AXILiteS_s_axi_U/n676 ,
         \Decision_AXILiteS_s_axi_U/n675 , \Decision_AXILiteS_s_axi_U/n674 ,
         \Decision_AXILiteS_s_axi_U/n673 , \Decision_AXILiteS_s_axi_U/n672 ,
         \Decision_AXILiteS_s_axi_U/n671 , \Decision_AXILiteS_s_axi_U/n670 ,
         \Decision_AXILiteS_s_axi_U/n669 , \Decision_AXILiteS_s_axi_U/n668 ,
         \Decision_AXILiteS_s_axi_U/n667 , \Decision_AXILiteS_s_axi_U/n666 ,
         \Decision_AXILiteS_s_axi_U/n665 , \Decision_AXILiteS_s_axi_U/n664 ,
         \Decision_AXILiteS_s_axi_U/n663 , \Decision_AXILiteS_s_axi_U/n662 ,
         \Decision_AXILiteS_s_axi_U/n661 , \Decision_AXILiteS_s_axi_U/n660 ,
         \Decision_AXILiteS_s_axi_U/n659 , \Decision_AXILiteS_s_axi_U/n658 ,
         \Decision_AXILiteS_s_axi_U/n657 , \Decision_AXILiteS_s_axi_U/n656 ,
         \Decision_AXILiteS_s_axi_U/n655 , \Decision_AXILiteS_s_axi_U/n654 ,
         \Decision_AXILiteS_s_axi_U/n653 , \Decision_AXILiteS_s_axi_U/n652 ,
         \Decision_AXILiteS_s_axi_U/n651 , \Decision_AXILiteS_s_axi_U/n650 ,
         \Decision_AXILiteS_s_axi_U/n649 , \Decision_AXILiteS_s_axi_U/n648 ,
         \Decision_AXILiteS_s_axi_U/n646 , \Decision_AXILiteS_s_axi_U/n645 ,
         \Decision_AXILiteS_s_axi_U/n644 , \Decision_AXILiteS_s_axi_U/n643 ,
         \Decision_AXILiteS_s_axi_U/n641 , \Decision_AXILiteS_s_axi_U/n640 ,
         \Decision_AXILiteS_s_axi_U/n639 , \Decision_AXILiteS_s_axi_U/n638 ,
         \Decision_AXILiteS_s_axi_U/n637 , \Decision_AXILiteS_s_axi_U/n636 ,
         \Decision_AXILiteS_s_axi_U/n635 , \Decision_AXILiteS_s_axi_U/n634 ,
         \Decision_AXILiteS_s_axi_U/n633 , \Decision_AXILiteS_s_axi_U/n632 ,
         \Decision_AXILiteS_s_axi_U/n631 , \Decision_AXILiteS_s_axi_U/n630 ,
         \Decision_AXILiteS_s_axi_U/n629 , \Decision_AXILiteS_s_axi_U/n628 ,
         \Decision_AXILiteS_s_axi_U/n627 , \Decision_AXILiteS_s_axi_U/n626 ,
         \Decision_AXILiteS_s_axi_U/n625 , \Decision_AXILiteS_s_axi_U/n624 ,
         \Decision_AXILiteS_s_axi_U/n623 , \Decision_AXILiteS_s_axi_U/n622 ,
         \Decision_AXILiteS_s_axi_U/n621 , \Decision_AXILiteS_s_axi_U/n620 ,
         \Decision_AXILiteS_s_axi_U/n619 , \Decision_AXILiteS_s_axi_U/n618 ,
         \Decision_AXILiteS_s_axi_U/n617 , \Decision_AXILiteS_s_axi_U/n616 ,
         \Decision_AXILiteS_s_axi_U/n615 , \Decision_AXILiteS_s_axi_U/n614 ,
         \Decision_AXILiteS_s_axi_U/n613 , \Decision_AXILiteS_s_axi_U/n612 ,
         \Decision_AXILiteS_s_axi_U/n611 , \Decision_AXILiteS_s_axi_U/n610 ,
         \Decision_AXILiteS_s_axi_U/n609 , \Decision_AXILiteS_s_axi_U/n608 ,
         \Decision_AXILiteS_s_axi_U/n607 , \Decision_AXILiteS_s_axi_U/n606 ,
         \Decision_AXILiteS_s_axi_U/n605 , \Decision_AXILiteS_s_axi_U/n604 ,
         \Decision_AXILiteS_s_axi_U/n603 , \Decision_AXILiteS_s_axi_U/n602 ,
         \Decision_AXILiteS_s_axi_U/n601 , \Decision_AXILiteS_s_axi_U/n600 ,
         \Decision_AXILiteS_s_axi_U/n599 , \Decision_AXILiteS_s_axi_U/n598 ,
         \Decision_AXILiteS_s_axi_U/n597 , \Decision_AXILiteS_s_axi_U/n596 ,
         \Decision_AXILiteS_s_axi_U/n595 , \Decision_AXILiteS_s_axi_U/n594 ,
         \Decision_AXILiteS_s_axi_U/n590 , \Decision_AXILiteS_s_axi_U/n586 ,
         \Decision_AXILiteS_s_axi_U/n582 , \Decision_AXILiteS_s_axi_U/n579 ,
         \Decision_AXILiteS_s_axi_U/n576 , \Decision_AXILiteS_s_axi_U/n575 ,
         \Decision_AXILiteS_s_axi_U/n574 , \Decision_AXILiteS_s_axi_U/n573 ,
         \Decision_AXILiteS_s_axi_U/n572 , \Decision_AXILiteS_s_axi_U/n571 ,
         \Decision_AXILiteS_s_axi_U/n570 , \Decision_AXILiteS_s_axi_U/n569 ,
         \Decision_AXILiteS_s_axi_U/n568 , \Decision_AXILiteS_s_axi_U/n567 ,
         \Decision_AXILiteS_s_axi_U/n566 , \Decision_AXILiteS_s_axi_U/n565 ,
         \Decision_AXILiteS_s_axi_U/n564 , \Decision_AXILiteS_s_axi_U/n563 ,
         \Decision_AXILiteS_s_axi_U/n562 , \Decision_AXILiteS_s_axi_U/n561 ,
         \Decision_AXILiteS_s_axi_U/n560 , \Decision_AXILiteS_s_axi_U/n559 ,
         \Decision_AXILiteS_s_axi_U/n558 , \Decision_AXILiteS_s_axi_U/n557 ,
         \Decision_AXILiteS_s_axi_U/n556 , \Decision_AXILiteS_s_axi_U/n555 ,
         \Decision_AXILiteS_s_axi_U/n554 , \Decision_AXILiteS_s_axi_U/n553 ,
         \Decision_AXILiteS_s_axi_U/n552 , \Decision_AXILiteS_s_axi_U/n551 ,
         \Decision_AXILiteS_s_axi_U/n550 , \Decision_AXILiteS_s_axi_U/n549 ,
         \Decision_AXILiteS_s_axi_U/n548 , \Decision_AXILiteS_s_axi_U/n547 ,
         \Decision_AXILiteS_s_axi_U/n546 , \Decision_AXILiteS_s_axi_U/n545 ,
         \Decision_AXILiteS_s_axi_U/n544 , \Decision_AXILiteS_s_axi_U/n543 ,
         \Decision_AXILiteS_s_axi_U/n542 , \Decision_AXILiteS_s_axi_U/n541 ,
         \Decision_AXILiteS_s_axi_U/n540 , \Decision_AXILiteS_s_axi_U/n539 ,
         \Decision_AXILiteS_s_axi_U/n538 , \Decision_AXILiteS_s_axi_U/n537 ,
         \Decision_AXILiteS_s_axi_U/n536 , \Decision_AXILiteS_s_axi_U/n535 ,
         \Decision_AXILiteS_s_axi_U/n533 , \Decision_AXILiteS_s_axi_U/n532 ,
         \Decision_AXILiteS_s_axi_U/n531 , \Decision_AXILiteS_s_axi_U/n530 ,
         \Decision_AXILiteS_s_axi_U/n529 , \Decision_AXILiteS_s_axi_U/n528 ,
         \Decision_AXILiteS_s_axi_U/n527 , \Decision_AXILiteS_s_axi_U/n526 ,
         \Decision_AXILiteS_s_axi_U/n525 , \Decision_AXILiteS_s_axi_U/n524 ,
         \Decision_AXILiteS_s_axi_U/n523 , \Decision_AXILiteS_s_axi_U/n522 ,
         \Decision_AXILiteS_s_axi_U/n521 , \Decision_AXILiteS_s_axi_U/n520 ,
         \Decision_AXILiteS_s_axi_U/n519 , \Decision_AXILiteS_s_axi_U/n518 ,
         \Decision_AXILiteS_s_axi_U/n517 , \Decision_AXILiteS_s_axi_U/n516 ,
         \Decision_AXILiteS_s_axi_U/n515 , \Decision_AXILiteS_s_axi_U/n514 ,
         \Decision_AXILiteS_s_axi_U/n513 , \Decision_AXILiteS_s_axi_U/n512 ,
         \Decision_AXILiteS_s_axi_U/n511 , \Decision_AXILiteS_s_axi_U/n510 ,
         \Decision_AXILiteS_s_axi_U/n509 , \Decision_AXILiteS_s_axi_U/n508 ,
         \Decision_AXILiteS_s_axi_U/n507 , \Decision_AXILiteS_s_axi_U/n506 ,
         \Decision_AXILiteS_s_axi_U/n505 , \Decision_AXILiteS_s_axi_U/n504 ,
         \Decision_AXILiteS_s_axi_U/n503 , \Decision_AXILiteS_s_axi_U/n502 ,
         \Decision_AXILiteS_s_axi_U/n501 , \Decision_AXILiteS_s_axi_U/n500 ,
         \Decision_AXILiteS_s_axi_U/n499 , \Decision_AXILiteS_s_axi_U/n498 ,
         \Decision_AXILiteS_s_axi_U/n497 , \Decision_AXILiteS_s_axi_U/n496 ,
         \Decision_AXILiteS_s_axi_U/n495 , \Decision_AXILiteS_s_axi_U/n494 ,
         \Decision_AXILiteS_s_axi_U/n493 , \Decision_AXILiteS_s_axi_U/n492 ,
         \Decision_AXILiteS_s_axi_U/n491 , \Decision_AXILiteS_s_axi_U/n490 ,
         \Decision_AXILiteS_s_axi_U/n489 , \Decision_AXILiteS_s_axi_U/n488 ,
         \Decision_AXILiteS_s_axi_U/n487 , \Decision_AXILiteS_s_axi_U/n486 ,
         \Decision_AXILiteS_s_axi_U/n485 , \Decision_AXILiteS_s_axi_U/n484 ,
         \Decision_AXILiteS_s_axi_U/n483 , \Decision_AXILiteS_s_axi_U/n482 ,
         \Decision_AXILiteS_s_axi_U/n481 , \Decision_AXILiteS_s_axi_U/n480 ,
         \Decision_AXILiteS_s_axi_U/n479 , \Decision_AXILiteS_s_axi_U/n478 ,
         \Decision_AXILiteS_s_axi_U/n477 , \Decision_AXILiteS_s_axi_U/n476 ,
         \Decision_AXILiteS_s_axi_U/n475 , \Decision_AXILiteS_s_axi_U/n474 ,
         \Decision_AXILiteS_s_axi_U/n473 , \Decision_AXILiteS_s_axi_U/n472 ,
         \Decision_AXILiteS_s_axi_U/n471 , \Decision_AXILiteS_s_axi_U/n470 ,
         \Decision_AXILiteS_s_axi_U/n469 , \Decision_AXILiteS_s_axi_U/n468 ,
         \Decision_AXILiteS_s_axi_U/n467 , \Decision_AXILiteS_s_axi_U/n466 ,
         \Decision_AXILiteS_s_axi_U/n465 , \Decision_AXILiteS_s_axi_U/n464 ,
         \Decision_AXILiteS_s_axi_U/n463 , \Decision_AXILiteS_s_axi_U/n462 ,
         \Decision_AXILiteS_s_axi_U/n461 , \Decision_AXILiteS_s_axi_U/n460 ,
         \Decision_AXILiteS_s_axi_U/n459 , \Decision_AXILiteS_s_axi_U/n458 ,
         \Decision_AXILiteS_s_axi_U/n457 , \Decision_AXILiteS_s_axi_U/n456 ,
         \Decision_AXILiteS_s_axi_U/n455 , \Decision_AXILiteS_s_axi_U/n454 ,
         \Decision_AXILiteS_s_axi_U/n453 , \Decision_AXILiteS_s_axi_U/n452 ,
         \Decision_AXILiteS_s_axi_U/n451 , \Decision_AXILiteS_s_axi_U/n450 ,
         \Decision_AXILiteS_s_axi_U/n449 , \Decision_AXILiteS_s_axi_U/n448 ,
         \Decision_AXILiteS_s_axi_U/n447 , \Decision_AXILiteS_s_axi_U/n446 ,
         \Decision_AXILiteS_s_axi_U/n445 , \Decision_AXILiteS_s_axi_U/n444 ,
         \Decision_AXILiteS_s_axi_U/n443 , \Decision_AXILiteS_s_axi_U/n442 ,
         \Decision_AXILiteS_s_axi_U/n441 , \Decision_AXILiteS_s_axi_U/n440 ,
         \Decision_AXILiteS_s_axi_U/n439 , \Decision_AXILiteS_s_axi_U/n438 ,
         \Decision_AXILiteS_s_axi_U/n437 , \Decision_AXILiteS_s_axi_U/n436 ,
         \Decision_AXILiteS_s_axi_U/n435 , \Decision_AXILiteS_s_axi_U/n434 ,
         \Decision_AXILiteS_s_axi_U/n433 , \Decision_AXILiteS_s_axi_U/n432 ,
         \Decision_AXILiteS_s_axi_U/n431 , \Decision_AXILiteS_s_axi_U/n430 ,
         \Decision_AXILiteS_s_axi_U/n429 , \Decision_AXILiteS_s_axi_U/n428 ,
         \Decision_AXILiteS_s_axi_U/n427 , \Decision_AXILiteS_s_axi_U/n426 ,
         \Decision_AXILiteS_s_axi_U/n425 , \Decision_AXILiteS_s_axi_U/n424 ,
         \Decision_AXILiteS_s_axi_U/n423 , \Decision_AXILiteS_s_axi_U/n422 ,
         \Decision_AXILiteS_s_axi_U/n421 , \Decision_AXILiteS_s_axi_U/n420 ,
         \Decision_AXILiteS_s_axi_U/n419 , \Decision_AXILiteS_s_axi_U/n418 ,
         \Decision_AXILiteS_s_axi_U/n417 , \Decision_AXILiteS_s_axi_U/n416 ,
         \Decision_AXILiteS_s_axi_U/n415 , \Decision_AXILiteS_s_axi_U/n414 ,
         \Decision_AXILiteS_s_axi_U/n413 , \Decision_AXILiteS_s_axi_U/n412 ,
         \Decision_AXILiteS_s_axi_U/n411 , \Decision_AXILiteS_s_axi_U/n410 ,
         \Decision_AXILiteS_s_axi_U/n409 , \Decision_AXILiteS_s_axi_U/n408 ,
         \Decision_AXILiteS_s_axi_U/n407 , \Decision_AXILiteS_s_axi_U/n406 ,
         \Decision_AXILiteS_s_axi_U/n405 , \Decision_AXILiteS_s_axi_U/n404 ,
         \Decision_AXILiteS_s_axi_U/n403 , \Decision_AXILiteS_s_axi_U/n402 ,
         \Decision_AXILiteS_s_axi_U/n401 , \Decision_AXILiteS_s_axi_U/n400 ,
         \Decision_AXILiteS_s_axi_U/n399 , \Decision_AXILiteS_s_axi_U/n398 ,
         \Decision_AXILiteS_s_axi_U/n397 , \Decision_AXILiteS_s_axi_U/n396 ,
         \Decision_AXILiteS_s_axi_U/n395 , \Decision_AXILiteS_s_axi_U/n394 ,
         \Decision_AXILiteS_s_axi_U/n393 , \Decision_AXILiteS_s_axi_U/n392 ,
         \Decision_AXILiteS_s_axi_U/n391 , \Decision_AXILiteS_s_axi_U/n390 ,
         \Decision_AXILiteS_s_axi_U/n389 , \Decision_AXILiteS_s_axi_U/n388 ,
         \Decision_AXILiteS_s_axi_U/n387 , \Decision_AXILiteS_s_axi_U/n386 ,
         \Decision_AXILiteS_s_axi_U/n385 , \Decision_AXILiteS_s_axi_U/n384 ,
         \Decision_AXILiteS_s_axi_U/n383 , \Decision_AXILiteS_s_axi_U/n382 ,
         \Decision_AXILiteS_s_axi_U/n381 , \Decision_AXILiteS_s_axi_U/n380 ,
         \Decision_AXILiteS_s_axi_U/n379 , \Decision_AXILiteS_s_axi_U/n378 ,
         \Decision_AXILiteS_s_axi_U/n377 , \Decision_AXILiteS_s_axi_U/n376 ,
         \Decision_AXILiteS_s_axi_U/n375 , \Decision_AXILiteS_s_axi_U/n374 ,
         \Decision_AXILiteS_s_axi_U/n373 , \Decision_AXILiteS_s_axi_U/n372 ,
         \Decision_AXILiteS_s_axi_U/n371 , \Decision_AXILiteS_s_axi_U/n370 ,
         \Decision_AXILiteS_s_axi_U/n369 , \Decision_AXILiteS_s_axi_U/n368 ,
         \Decision_AXILiteS_s_axi_U/n367 , \Decision_AXILiteS_s_axi_U/n366 ,
         \Decision_AXILiteS_s_axi_U/n365 , \Decision_AXILiteS_s_axi_U/n364 ,
         \Decision_AXILiteS_s_axi_U/n363 , \Decision_AXILiteS_s_axi_U/n362 ,
         \Decision_AXILiteS_s_axi_U/n361 , \Decision_AXILiteS_s_axi_U/n360 ,
         \Decision_AXILiteS_s_axi_U/n359 , \Decision_AXILiteS_s_axi_U/n358 ,
         \Decision_AXILiteS_s_axi_U/n357 , \Decision_AXILiteS_s_axi_U/n356 ,
         \Decision_AXILiteS_s_axi_U/n355 , \Decision_AXILiteS_s_axi_U/n354 ,
         \Decision_AXILiteS_s_axi_U/n353 , \Decision_AXILiteS_s_axi_U/n352 ,
         \Decision_AXILiteS_s_axi_U/n351 , \Decision_AXILiteS_s_axi_U/n350 ,
         \Decision_AXILiteS_s_axi_U/n349 , \Decision_AXILiteS_s_axi_U/n348 ,
         \Decision_AXILiteS_s_axi_U/n347 , \Decision_AXILiteS_s_axi_U/n346 ,
         \Decision_AXILiteS_s_axi_U/n345 , \Decision_AXILiteS_s_axi_U/n344 ,
         \Decision_AXILiteS_s_axi_U/n343 , \Decision_AXILiteS_s_axi_U/n342 ,
         \Decision_AXILiteS_s_axi_U/n341 , \Decision_AXILiteS_s_axi_U/n340 ,
         \Decision_AXILiteS_s_axi_U/n339 , \Decision_AXILiteS_s_axi_U/n338 ,
         \Decision_AXILiteS_s_axi_U/n337 , \Decision_AXILiteS_s_axi_U/n336 ,
         \Decision_AXILiteS_s_axi_U/n335 , \Decision_AXILiteS_s_axi_U/n334 ,
         \Decision_AXILiteS_s_axi_U/n333 , \Decision_AXILiteS_s_axi_U/n332 ,
         \Decision_AXILiteS_s_axi_U/n331 , \Decision_AXILiteS_s_axi_U/n330 ,
         \Decision_AXILiteS_s_axi_U/n329 , \Decision_AXILiteS_s_axi_U/n328 ,
         \Decision_AXILiteS_s_axi_U/n327 , \Decision_AXILiteS_s_axi_U/n326 ,
         \Decision_AXILiteS_s_axi_U/n325 , \Decision_AXILiteS_s_axi_U/n324 ,
         \Decision_AXILiteS_s_axi_U/n323 , \Decision_AXILiteS_s_axi_U/n322 ,
         \Decision_AXILiteS_s_axi_U/n321 , \Decision_AXILiteS_s_axi_U/n320 ,
         \Decision_AXILiteS_s_axi_U/n319 , \Decision_AXILiteS_s_axi_U/n318 ,
         \Decision_AXILiteS_s_axi_U/n317 , \Decision_AXILiteS_s_axi_U/n316 ,
         \Decision_AXILiteS_s_axi_U/n315 , \Decision_AXILiteS_s_axi_U/n313 ,
         \Decision_AXILiteS_s_axi_U/n312 , \Decision_AXILiteS_s_axi_U/n311 ,
         \Decision_AXILiteS_s_axi_U/n310 , \Decision_AXILiteS_s_axi_U/n309 ,
         \Decision_AXILiteS_s_axi_U/n308 , \Decision_AXILiteS_s_axi_U/n307 ,
         \Decision_AXILiteS_s_axi_U/n306 , \Decision_AXILiteS_s_axi_U/n305 ,
         \Decision_AXILiteS_s_axi_U/n304 , \Decision_AXILiteS_s_axi_U/n303 ,
         \Decision_AXILiteS_s_axi_U/n302 , \Decision_AXILiteS_s_axi_U/n301 ,
         \Decision_AXILiteS_s_axi_U/n299 , \Decision_AXILiteS_s_axi_U/n298 ,
         \Decision_AXILiteS_s_axi_U/n297 , \Decision_AXILiteS_s_axi_U/n296 ,
         \Decision_AXILiteS_s_axi_U/n295 , \Decision_AXILiteS_s_axi_U/n294 ,
         \Decision_AXILiteS_s_axi_U/n293 , \Decision_AXILiteS_s_axi_U/n292 ,
         \Decision_AXILiteS_s_axi_U/n291 , \Decision_AXILiteS_s_axi_U/n290 ,
         \Decision_AXILiteS_s_axi_U/n289 , \Decision_AXILiteS_s_axi_U/n288 ,
         \Decision_AXILiteS_s_axi_U/n287 , \Decision_AXILiteS_s_axi_U/n286 ,
         \Decision_AXILiteS_s_axi_U/n285 , \Decision_AXILiteS_s_axi_U/n284 ,
         \Decision_AXILiteS_s_axi_U/n283 , \Decision_AXILiteS_s_axi_U/n282 ,
         \Decision_AXILiteS_s_axi_U/n281 , \Decision_AXILiteS_s_axi_U/n280 ,
         \Decision_AXILiteS_s_axi_U/n279 , \Decision_AXILiteS_s_axi_U/n278 ,
         \Decision_AXILiteS_s_axi_U/n277 , \Decision_AXILiteS_s_axi_U/n276 ,
         \Decision_AXILiteS_s_axi_U/n275 , \Decision_AXILiteS_s_axi_U/n274 ,
         \Decision_AXILiteS_s_axi_U/n273 , \Decision_AXILiteS_s_axi_U/n272 ,
         \Decision_AXILiteS_s_axi_U/n271 , \Decision_AXILiteS_s_axi_U/n270 ,
         \Decision_AXILiteS_s_axi_U/n269 , \Decision_AXILiteS_s_axi_U/n268 ,
         \Decision_AXILiteS_s_axi_U/n267 , \Decision_AXILiteS_s_axi_U/n266 ,
         \Decision_AXILiteS_s_axi_U/n265 , \Decision_AXILiteS_s_axi_U/n264 ,
         \Decision_AXILiteS_s_axi_U/n263 , \Decision_AXILiteS_s_axi_U/n262 ,
         \Decision_AXILiteS_s_axi_U/n261 , \Decision_AXILiteS_s_axi_U/n260 ,
         \Decision_AXILiteS_s_axi_U/n259 , \Decision_AXILiteS_s_axi_U/n258 ,
         \Decision_AXILiteS_s_axi_U/n257 , \Decision_AXILiteS_s_axi_U/n256 ,
         \Decision_AXILiteS_s_axi_U/n255 , \Decision_AXILiteS_s_axi_U/n254 ,
         \Decision_AXILiteS_s_axi_U/n253 , \Decision_AXILiteS_s_axi_U/n252 ,
         \Decision_AXILiteS_s_axi_U/n251 , \Decision_AXILiteS_s_axi_U/n250 ,
         \Decision_AXILiteS_s_axi_U/n249 , \Decision_AXILiteS_s_axi_U/n248 ,
         \Decision_AXILiteS_s_axi_U/n247 , \Decision_AXILiteS_s_axi_U/n246 ,
         \Decision_AXILiteS_s_axi_U/n245 , \Decision_AXILiteS_s_axi_U/n244 ,
         \Decision_AXILiteS_s_axi_U/n243 , \Decision_AXILiteS_s_axi_U/n242 ,
         \Decision_AXILiteS_s_axi_U/n241 , \Decision_AXILiteS_s_axi_U/n240 ,
         \Decision_AXILiteS_s_axi_U/n239 , \Decision_AXILiteS_s_axi_U/n238 ,
         \Decision_AXILiteS_s_axi_U/n237 , \Decision_AXILiteS_s_axi_U/n236 ,
         \Decision_AXILiteS_s_axi_U/n235 , \Decision_AXILiteS_s_axi_U/n234 ,
         \Decision_AXILiteS_s_axi_U/n233 , \Decision_AXILiteS_s_axi_U/n232 ,
         \Decision_AXILiteS_s_axi_U/n231 , \Decision_AXILiteS_s_axi_U/n230 ,
         \Decision_AXILiteS_s_axi_U/n229 , \Decision_AXILiteS_s_axi_U/n228 ,
         \Decision_AXILiteS_s_axi_U/n227 , \Decision_AXILiteS_s_axi_U/n226 ,
         \Decision_AXILiteS_s_axi_U/n225 , \Decision_AXILiteS_s_axi_U/n224 ,
         \Decision_AXILiteS_s_axi_U/n223 , \Decision_AXILiteS_s_axi_U/n222 ,
         \Decision_AXILiteS_s_axi_U/n221 , \Decision_AXILiteS_s_axi_U/n220 ,
         \Decision_AXILiteS_s_axi_U/n219 , \Decision_AXILiteS_s_axi_U/n218 ,
         \Decision_AXILiteS_s_axi_U/n217 , \Decision_AXILiteS_s_axi_U/n216 ,
         \Decision_AXILiteS_s_axi_U/n215 , \Decision_AXILiteS_s_axi_U/n214 ,
         \Decision_AXILiteS_s_axi_U/n213 , \Decision_AXILiteS_s_axi_U/n212 ,
         \Decision_AXILiteS_s_axi_U/n211 , \Decision_AXILiteS_s_axi_U/n210 ,
         \Decision_AXILiteS_s_axi_U/n209 , \Decision_AXILiteS_s_axi_U/n208 ,
         \Decision_AXILiteS_s_axi_U/n207 , \Decision_AXILiteS_s_axi_U/n206 ,
         \Decision_AXILiteS_s_axi_U/n205 , \Decision_AXILiteS_s_axi_U/n204 ,
         \Decision_AXILiteS_s_axi_U/n203 , \Decision_AXILiteS_s_axi_U/n202 ,
         \Decision_AXILiteS_s_axi_U/n201 , \Decision_AXILiteS_s_axi_U/n200 ,
         \Decision_AXILiteS_s_axi_U/n199 , \Decision_AXILiteS_s_axi_U/n198 ,
         \Decision_AXILiteS_s_axi_U/n197 , \Decision_AXILiteS_s_axi_U/n196 ,
         \Decision_AXILiteS_s_axi_U/n195 , \Decision_AXILiteS_s_axi_U/n194 ,
         \Decision_AXILiteS_s_axi_U/n193 , \Decision_AXILiteS_s_axi_U/n192 ,
         \Decision_AXILiteS_s_axi_U/n191 , \Decision_AXILiteS_s_axi_U/n190 ,
         \Decision_AXILiteS_s_axi_U/n189 , \Decision_AXILiteS_s_axi_U/n188 ,
         \Decision_AXILiteS_s_axi_U/n187 , \Decision_AXILiteS_s_axi_U/n186 ,
         \Decision_AXILiteS_s_axi_U/n185 , \Decision_AXILiteS_s_axi_U/n184 ,
         \Decision_AXILiteS_s_axi_U/n183 , \Decision_AXILiteS_s_axi_U/n182 ,
         \Decision_AXILiteS_s_axi_U/n181 , \Decision_AXILiteS_s_axi_U/n180 ,
         \Decision_AXILiteS_s_axi_U/n179 , \Decision_AXILiteS_s_axi_U/n178 ,
         \Decision_AXILiteS_s_axi_U/n177 , \Decision_AXILiteS_s_axi_U/n176 ,
         \Decision_AXILiteS_s_axi_U/n175 , \Decision_AXILiteS_s_axi_U/n174 ,
         \Decision_AXILiteS_s_axi_U/n173 , \Decision_AXILiteS_s_axi_U/n172 ,
         \Decision_AXILiteS_s_axi_U/n171 , \Decision_AXILiteS_s_axi_U/n170 ,
         \Decision_AXILiteS_s_axi_U/n169 , \Decision_AXILiteS_s_axi_U/n168 ,
         \Decision_AXILiteS_s_axi_U/n167 , \Decision_AXILiteS_s_axi_U/n166 ,
         \Decision_AXILiteS_s_axi_U/n165 , \Decision_AXILiteS_s_axi_U/n164 ,
         \Decision_AXILiteS_s_axi_U/n163 , \Decision_AXILiteS_s_axi_U/n162 ,
         \Decision_AXILiteS_s_axi_U/n161 , \Decision_AXILiteS_s_axi_U/n160 ,
         \Decision_AXILiteS_s_axi_U/n159 , \Decision_AXILiteS_s_axi_U/n158 ,
         \Decision_AXILiteS_s_axi_U/n157 , \Decision_AXILiteS_s_axi_U/n155 ,
         \Decision_AXILiteS_s_axi_U/n154 , \Decision_AXILiteS_s_axi_U/n153 ,
         \Decision_AXILiteS_s_axi_U/n152 ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[0] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[1] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[2] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[3] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[4] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[5] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[6] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[7] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[8] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[9] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[10] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[11] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[12] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[13] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[14] ,
         \Decision_AXILiteS_s_axi_U/int_ap_return[15] ,
         \Decision_AXILiteS_s_axi_U/int_isr[0] ,
         \Decision_AXILiteS_s_axi_U/int_isr[1] ,
         \Decision_AXILiteS_s_axi_U/int_ier[0] ,
         \Decision_AXILiteS_s_axi_U/int_ier[1] ,
         \Decision_AXILiteS_s_axi_U/int_gie ,
         \Decision_AXILiteS_s_axi_U/int_auto_restart ,
         \Decision_AXILiteS_s_axi_U/int_ap_done ,
         \Decision_AXILiteS_s_axi_U/rstate[0] ,
         \Decision_AXILiteS_s_axi_U/waddr[0] ,
         \Decision_AXILiteS_s_axi_U/waddr[1] ,
         \Decision_AXILiteS_s_axi_U/waddr[2] ,
         \Decision_AXILiteS_s_axi_U/waddr[3] ,
         \Decision_AXILiteS_s_axi_U/waddr[4] ,
         \Decision_AXILiteS_s_axi_U/waddr[5] ,
         \Decision_AXILiteS_s_axi_U/waddr[6] ,
         \Decision_AXILiteS_s_axi_U/wstate[0] ,
         \Decision_AXILiteS_s_axi_U/wstate[1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1228 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1227 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1226 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1225 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1224 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1223 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1222 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1221 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1220 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1219 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1218 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1217 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1216 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1215 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1214 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1213 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1212 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1211 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1210 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1209 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1208 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1207 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1206 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1205 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1204 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1203 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1202 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1201 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1200 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1199 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1198 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1197 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1196 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1195 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1194 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1193 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1192 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1191 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1190 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1189 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1188 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1187 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1186 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1185 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1184 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1183 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1182 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1181 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1180 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1179 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1178 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1177 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1176 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1175 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1174 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1173 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1172 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1171 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1170 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1169 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1168 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1167 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1166 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1165 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1164 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1163 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1162 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1161 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1160 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1159 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1158 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1157 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1156 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1155 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1154 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1153 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1152 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1151 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1150 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1149 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1148 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1147 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1146 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1145 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1144 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1143 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1142 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1141 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1140 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1139 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1138 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1137 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1136 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1135 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1134 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1133 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1132 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1131 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1130 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1129 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1128 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1127 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1126 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1125 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1124 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1123 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1122 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1121 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1120 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1119 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1118 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1117 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1116 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1115 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1114 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1113 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1112 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1111 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1110 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1109 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1108 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1107 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1106 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1105 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1104 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1103 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1102 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1101 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1100 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1099 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1098 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1097 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1096 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1095 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1094 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1093 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1092 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1091 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1090 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1089 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1088 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1087 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1086 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1085 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1084 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1083 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1082 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1081 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1080 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1079 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1078 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1077 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1076 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1075 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1074 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1073 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1072 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1071 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1070 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1069 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1068 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1067 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1066 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1065 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1064 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1063 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1062 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1061 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1060 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1059 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1058 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1057 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1056 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1055 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1054 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1053 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1052 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1051 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1050 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1049 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1048 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1047 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1046 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1045 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1044 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1043 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1042 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1041 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1040 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1039 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1038 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1037 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1036 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1035 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1034 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1033 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1032 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1031 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1030 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1029 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1028 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1027 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1026 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1025 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1024 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1023 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1022 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1021 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1020 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1019 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1018 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1017 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1016 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1015 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1014 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1013 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1012 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1011 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1010 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1009 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1008 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1007 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1006 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1005 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1004 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1003 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1002 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1001 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1000 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n999 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n998 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n997 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n996 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n995 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n994 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n993 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n992 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n991 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n990 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n989 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n988 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n987 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n986 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n985 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n984 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n983 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n982 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n981 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n980 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n979 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n978 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n977 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n976 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n975 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n974 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n973 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n972 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n971 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n970 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n969 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n968 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n967 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n966 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n965 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n964 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n963 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n962 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n961 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n960 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n959 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n958 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n957 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n956 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n955 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n954 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n953 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n952 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n951 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n950 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n949 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n948 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n947 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n946 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n945 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n944 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n943 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n942 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n941 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n940 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n939 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n938 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n937 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n936 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n935 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n934 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n933 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n932 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n931 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n930 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n929 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n928 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n927 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n926 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n925 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n924 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n923 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n922 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n921 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n920 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n919 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n918 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n917 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n916 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n915 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n914 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n913 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n912 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n911 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n910 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n909 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n908 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n907 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n906 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n905 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n904 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n903 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n902 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n901 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n900 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n899 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n898 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n897 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n896 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n895 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n894 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n893 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n892 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n890 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n888 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n886 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n884 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n882 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n880 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n878 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n876 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n874 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n872 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n870 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n868 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n866 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n864 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n862 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n859 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n858 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n857 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n856 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n855 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n854 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n853 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n852 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n851 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n850 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n849 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n848 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n847 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n846 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n845 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n844 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n842 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n841 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n840 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n839 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n838 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n837 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n836 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n835 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n834 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n833 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n832 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n831 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n830 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n829 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n828 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n827 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n825 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n824 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n823 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n822 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n821 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n820 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n819 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n818 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n817 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n816 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n815 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n814 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n813 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n812 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n811 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n810 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n809 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n807 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n806 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n804 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n802 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n800 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n798 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n796 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n794 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n792 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n790 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n788 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n786 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n784 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n782 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n780 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n778 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n776 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n773 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n772 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n771 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n770 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n769 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n768 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n767 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n766 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n765 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n764 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n763 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n762 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n761 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n760 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n759 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n758 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n757 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n756 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n755 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n754 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n753 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n752 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n751 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n750 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n749 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n748 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n747 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n746 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n745 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n744 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n743 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n742 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n741 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n740 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n739 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n738 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n737 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n736 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n735 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n734 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n733 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n732 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n731 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n730 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n729 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n728 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n727 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n726 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n725 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n724 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n723 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n722 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n721 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n720 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n719 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n718 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n717 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n716 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n715 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n714 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n713 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n712 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n711 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n710 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n709 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n708 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n707 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n706 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n705 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n704 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n703 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n702 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n701 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n700 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n699 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n698 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n697 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n696 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n695 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n694 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n693 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n692 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n691 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n690 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n689 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n688 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n687 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n686 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n685 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n684 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n683 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n682 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n681 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n680 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n679 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n678 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n677 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n676 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n675 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n674 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n673 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n672 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n671 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n670 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n669 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n668 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n667 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n666 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n665 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n664 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n663 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n662 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n661 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n660 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n659 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n658 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n657 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n656 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n655 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n654 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n653 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n652 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n650 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n649 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n648 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n646 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n644 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n642 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n640 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n638 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n636 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n634 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n632 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n630 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n628 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n626 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n624 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n622 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n620 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n618 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n615 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n614 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n612 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n610 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n608 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n606 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n604 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n602 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n600 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n598 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n596 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n594 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n592 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n590 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n588 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n586 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n584 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n581 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n579 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n577 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n575 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n573 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n571 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n569 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n567 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n565 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n563 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n561 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n559 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n557 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n555 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n553 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n551 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n550 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n547 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n546 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n544 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n542 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n540 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n538 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n536 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n534 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n532 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n530 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n528 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n526 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n524 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n522 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n520 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n518 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n516 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n513 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n512 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n510 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n508 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n506 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n504 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n502 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n500 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n498 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n496 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n494 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n492 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n490 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n488 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n486 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n484 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n482 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n479 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n478 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n476 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n474 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n472 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n470 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n468 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n466 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n464 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n462 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n460 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n458 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n456 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n454 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n452 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n450 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n448 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n445 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n444 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n442 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n440 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n438 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n436 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n434 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n432 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n430 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n428 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n426 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n424 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n422 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n420 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n418 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n416 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n414 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n411 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n410 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n409 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n407 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n405 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n403 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n401 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n399 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n397 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n395 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n393 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n391 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n389 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n387 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n385 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n383 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n381 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n379 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n375 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n373 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n372 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n371 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n370 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n369 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n368 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n367 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n365 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n363 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n362 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n361 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n359 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n358 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n357 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n356 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n355 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n354 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n352 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n351 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n350 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n349 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n348 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n347 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n346 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n345 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n344 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n343 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n342 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n341 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n340 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n339 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n338 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n337 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n336 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n335 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n334 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n333 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n332 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n331 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n330 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n329 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n328 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n327 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n326 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n325 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n324 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n323 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n322 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n321 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n320 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n319 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n318 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n317 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n316 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n315 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n314 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n313 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n312 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n311 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n310 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n309 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n308 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n307 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n306 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n305 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n304 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n303 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n302 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n301 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n300 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n299 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n298 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n297 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n296 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n295 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n294 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n293 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n292 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n291 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n290 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n289 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n288 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n287 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n286 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n285 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n284 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n283 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n282 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n281 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n280 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n279 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n278 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n277 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n276 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n275 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n274 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n273 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n272 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n271 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n270 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n269 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n268 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n267 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n266 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n265 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n264 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n263 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n262 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n261 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n260 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n259 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n258 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n257 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n256 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n255 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n254 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n253 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n252 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n251 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n250 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n249 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n248 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n247 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n246 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n245 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n244 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n243 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n242 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n241 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n240 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n239 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n238 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n237 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n236 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n235 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n234 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n233 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n232 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n231 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n230 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n229 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n228 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n227 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n226 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n225 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n224 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n223 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n222 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n221 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n220 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n219 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n218 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n217 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n216 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n215 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n214 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n213 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n212 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n211 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n210 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n209 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n208 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n207 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n206 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n205 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n204 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n203 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n202 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n201 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n200 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n199 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n198 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n197 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n196 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n195 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n194 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n193 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n192 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n191 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n190 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n189 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n188 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n187 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n186 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n185 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n184 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n183 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n182 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n181 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n180 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n179 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n178 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n177 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n176 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n175 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n174 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n173 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n172 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n171 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n170 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n169 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n168 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n167 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n166 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n165 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n164 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n163 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n162 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n161 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n160 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n159 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n158 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n157 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n156 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n155 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n154 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n153 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n152 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n151 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n150 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n149 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n148 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n147 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n146 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n145 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n144 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n143 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n142 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n141 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n140 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n139 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n138 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n137 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n136 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n135 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n134 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n133 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n132 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n131 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n130 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n129 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n128 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n127 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n126 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n125 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n124 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n123 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n122 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n121 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n120 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n119 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n118 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n117 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n116 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n115 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n114 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n113 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n112 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n111 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n110 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n109 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n108 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n107 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n106 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n105 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n104 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n103 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n102 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n101 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n100 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n99 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n98 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n97 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n96 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n95 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n94 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n93 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n92 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n91 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n90 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n89 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n88 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n87 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n86 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n85 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n84 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n83 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n82 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n81 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n80 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n79 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n78 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n77 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n76 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n75 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n74 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n73 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n72 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n71 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n70 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n69 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n68 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n67 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n66 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n65 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n64 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n63 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n62 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n61 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n60 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n59 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n58 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n57 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n56 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n55 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n54 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n53 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n52 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n51 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n50 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n49 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n48 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n47 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n46 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n45 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n38 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n37 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n36 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n32 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n31 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n30 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n29 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n28 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n27 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n26 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n25 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n24 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n20 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n19 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n18 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n17 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n15 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n14 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n13 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n12 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n11 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n10 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n9 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n8 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n6 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n5 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n3 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n2 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1 ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][15] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][0] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][1] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][2] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][3] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][4] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][5] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][6] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][7] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][8] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][9] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][10] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][11] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][12] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][13] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][14] ,
         \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][15] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n162 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n161 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n160 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n159 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n158 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n157 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n156 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n155 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n154 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n153 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n152 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n151 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n150 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n149 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n148 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n147 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n146 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n145 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n144 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n143 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n142 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n141 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n140 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n139 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n138 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n137 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n136 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n135 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n134 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n133 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n132 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n131 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n130 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n129 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n128 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n127 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n126 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n125 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n124 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n123 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n122 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n121 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n120 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n119 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n118 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n117 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n116 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n115 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n114 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n113 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n112 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n111 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n110 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n109 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n108 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n107 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n106 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n105 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n104 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n103 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n102 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n101 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n100 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n99 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n98 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n97 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n96 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n95 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n94 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n93 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n92 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n91 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n90 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n89 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n88 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n87 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n86 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n85 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n83 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n82 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n81 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n80 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n79 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n76 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n75 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n73 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n71 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n70 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n69 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n68 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n67 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n66 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n65 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n64 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n63 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n62 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n60 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n59 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n58 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n57 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n56 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n55 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n54 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n53 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n52 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n51 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n49 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n48 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n47 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n46 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n45 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n44 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n43 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n42 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n41 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n40 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n39 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n38 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n37 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n36 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n35 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n34 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n33 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n32 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n31 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n30 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n29 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n26 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n25 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n24 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n23 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n21 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n20 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n19 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n18 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n16 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n15 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n14 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n13 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n12 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n9 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n8 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n7 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n6 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n4 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n3 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/n1 ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ,
         \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n162 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n161 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n160 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n159 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n158 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n157 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n156 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n155 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n154 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n153 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n152 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n151 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n150 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n149 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n148 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n147 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n146 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n145 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n144 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n143 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n142 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n141 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n140 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n139 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n138 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n137 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n136 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n135 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n134 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n133 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n132 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n131 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n130 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n129 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n128 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n127 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n126 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n125 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n124 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n123 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n122 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n121 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n120 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n119 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n118 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n117 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n116 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n115 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n114 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n113 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n112 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n111 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n110 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n109 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n108 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n107 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n106 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n105 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n104 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n103 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n102 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n101 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n100 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n99 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n98 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n97 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n96 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n95 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n94 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n93 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n92 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n91 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n90 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n89 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n88 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n87 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n85 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n84 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n83 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n82 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n81 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n78 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n77 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n75 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n73 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n72 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n71 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n70 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n69 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n68 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n67 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n66 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n65 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n64 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n62 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n61 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n60 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n59 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n58 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n57 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n56 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n55 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n54 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n53 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n51 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n50 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n49 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n48 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n47 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n46 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n45 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n44 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n43 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n42 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n41 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n40 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n39 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n38 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n37 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n36 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n35 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n34 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n32 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n31 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n30 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n29 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n27 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n26 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n25 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n24 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n22 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n21 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n20 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n19 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n17 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n16 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n15 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n13 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n12 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n11 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n9 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n8 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n7 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n6 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n4 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n3 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/n1 ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ,
         \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ,
         \dp_cluster_1/add_1107_aco/carry[31] ,
         \dp_cluster_1/add_1107_aco/carry[30] ,
         \dp_cluster_1/add_1107_aco/carry[29] ,
         \dp_cluster_1/add_1107_aco/carry[28] ,
         \dp_cluster_1/add_1107_aco/carry[27] ,
         \dp_cluster_1/add_1107_aco/carry[26] ,
         \dp_cluster_1/add_1107_aco/carry[25] ,
         \dp_cluster_1/add_1107_aco/carry[24] ,
         \dp_cluster_1/add_1107_aco/carry[23] ,
         \dp_cluster_1/add_1107_aco/carry[22] ,
         \dp_cluster_1/add_1107_aco/carry[21] ,
         \dp_cluster_1/add_1107_aco/carry[20] ,
         \dp_cluster_1/add_1107_aco/carry[19] ,
         \dp_cluster_1/add_1107_aco/carry[18] ,
         \dp_cluster_1/add_1107_aco/carry[17] ,
         \dp_cluster_1/add_1107_aco/carry[16] ,
         \dp_cluster_1/add_1107_aco/carry[15] ,
         \dp_cluster_1/add_1107_aco/carry[14] ,
         \dp_cluster_1/add_1107_aco/carry[13] ,
         \dp_cluster_1/add_1107_aco/carry[12] ,
         \dp_cluster_1/add_1107_aco/carry[11] ,
         \dp_cluster_1/add_1107_aco/carry[10] ,
         \dp_cluster_1/add_1107_aco/carry[9] ,
         \dp_cluster_1/add_1107_aco/carry[8] ,
         \dp_cluster_1/add_1107_aco/carry[7] ,
         \dp_cluster_1/add_1107_aco/carry[6] ,
         \dp_cluster_1/add_1107_aco/carry[5] ,
         \dp_cluster_1/add_1107_aco/carry[4] ,
         \dp_cluster_1/add_1107_aco/carry[3] ,
         \dp_cluster_1/add_1107_aco/carry[2] ,
         \dp_cluster_0/add_1147_aco/carry[31] ,
         \dp_cluster_0/add_1147_aco/carry[30] ,
         \dp_cluster_0/add_1147_aco/carry[29] ,
         \dp_cluster_0/add_1147_aco/carry[28] ,
         \dp_cluster_0/add_1147_aco/carry[27] ,
         \dp_cluster_0/add_1147_aco/carry[26] ,
         \dp_cluster_0/add_1147_aco/carry[25] ,
         \dp_cluster_0/add_1147_aco/carry[24] ,
         \dp_cluster_0/add_1147_aco/carry[23] ,
         \dp_cluster_0/add_1147_aco/carry[22] ,
         \dp_cluster_0/add_1147_aco/carry[21] ,
         \dp_cluster_0/add_1147_aco/carry[20] ,
         \dp_cluster_0/add_1147_aco/carry[19] ,
         \dp_cluster_0/add_1147_aco/carry[18] ,
         \dp_cluster_0/add_1147_aco/carry[17] ,
         \dp_cluster_0/add_1147_aco/carry[16] ,
         \dp_cluster_0/add_1147_aco/carry[15] ,
         \dp_cluster_0/add_1147_aco/carry[14] ,
         \dp_cluster_0/add_1147_aco/carry[13] ,
         \dp_cluster_0/add_1147_aco/carry[12] ,
         \dp_cluster_0/add_1147_aco/carry[11] ,
         \dp_cluster_0/add_1147_aco/carry[10] ,
         \dp_cluster_0/add_1147_aco/carry[9] ,
         \dp_cluster_0/add_1147_aco/carry[8] ,
         \dp_cluster_0/add_1147_aco/carry[7] ,
         \dp_cluster_0/add_1147_aco/carry[6] ,
         \dp_cluster_0/add_1147_aco/carry[5] ,
         \dp_cluster_0/add_1147_aco/carry[4] ,
         \dp_cluster_0/add_1147_aco/carry[3] ,
         \dp_cluster_0/add_1147_aco/carry[2] , \add_1415/carry[31] ,
         \add_1415/carry[30] , \add_1415/carry[29] , \add_1415/carry[28] ,
         \add_1415/carry[27] , \add_1415/carry[26] , \add_1415/carry[25] ,
         \add_1415/carry[24] , \add_1415/carry[23] , \add_1415/carry[22] ,
         \add_1415/carry[21] , \add_1415/carry[20] , \add_1415/carry[19] ,
         \add_1415/carry[18] , \add_1415/carry[17] , \add_1415/carry[16] ,
         \add_1415/carry[15] , \add_1415/carry[14] , \add_1415/carry[13] ,
         \add_1415/carry[12] , \add_1415/carry[11] , \add_1415/carry[10] ,
         \add_1415/carry[9] , \add_1415/carry[8] , \add_1415/carry[7] ,
         \add_1415/carry[6] , \add_1415/carry[5] , \add_1415/carry[4] ,
         \add_1415/carry[3] , \add_1415/carry[2] , \add_1413/carry[31] ,
         \add_1413/carry[30] , \add_1413/carry[29] , \add_1413/carry[28] ,
         \add_1413/carry[27] , \add_1413/carry[26] , \add_1413/carry[25] ,
         \add_1413/carry[24] , \add_1413/carry[23] , \add_1413/carry[22] ,
         \add_1413/carry[21] , \add_1413/carry[20] , \add_1413/carry[19] ,
         \add_1413/carry[18] , \add_1413/carry[17] , \add_1413/carry[16] ,
         \add_1413/carry[15] , \add_1413/carry[14] , \add_1413/carry[13] ,
         \add_1413/carry[12] , \add_1413/carry[11] , \add_1413/carry[10] ,
         \add_1413/carry[9] , \add_1413/carry[8] , \add_1413/carry[7] ,
         \add_1413/carry[6] , \add_1413/carry[5] , \add_1413/carry[4] ,
         \add_1413/carry[3] , \add_1413/carry[2] , \add_1407/carry[31] ,
         \add_1407/carry[30] , \add_1407/carry[29] , \add_1407/carry[28] ,
         \add_1407/carry[27] , \add_1407/carry[26] , \add_1407/carry[25] ,
         \add_1407/carry[24] , \add_1407/carry[23] , \add_1407/carry[22] ,
         \add_1407/carry[21] , \add_1407/carry[20] , \add_1407/carry[19] ,
         \add_1407/carry[18] , \add_1407/carry[17] , \add_1407/carry[16] ,
         \add_1407/carry[15] , \add_1407/carry[14] , \add_1407/carry[13] ,
         \add_1407/carry[12] , \add_1407/carry[11] , \add_1407/carry[10] ,
         \add_1407/carry[9] , \add_1407/carry[8] , \add_1407/carry[7] ,
         \add_1407/carry[6] , \add_1407/carry[5] , \add_1407/carry[4] ,
         \add_1407/carry[3] , \add_1407/carry[2] , \add_1405/carry[31] ,
         \add_1405/carry[30] , \add_1405/carry[29] , \add_1405/carry[28] ,
         \add_1405/carry[27] , \add_1405/carry[26] , \add_1405/carry[25] ,
         \add_1405/carry[24] , \add_1405/carry[23] , \add_1405/carry[22] ,
         \add_1405/carry[21] , \add_1405/carry[20] , \add_1405/carry[19] ,
         \add_1405/carry[18] , \add_1405/carry[17] , \add_1405/carry[16] ,
         \add_1405/carry[15] , \add_1405/carry[14] , \add_1405/carry[13] ,
         \add_1405/carry[12] , \add_1405/carry[11] , \add_1405/carry[10] ,
         \add_1405/carry[9] , \add_1405/carry[8] , \add_1405/carry[7] ,
         \add_1405/carry[6] , \add_1405/carry[5] , \add_1405/carry[4] ,
         \add_1405/carry[3] , \add_1405/carry[2] , \add_1393/carry[31] ,
         \add_1393/carry[30] , \add_1393/carry[29] , \add_1393/carry[28] ,
         \add_1393/carry[27] , \add_1393/carry[26] , \add_1393/carry[25] ,
         \add_1393/carry[24] , \add_1393/carry[23] , \add_1393/carry[22] ,
         \add_1393/carry[21] , \add_1393/carry[20] , \add_1393/carry[19] ,
         \add_1393/carry[18] , \add_1393/carry[17] , \add_1393/carry[16] ,
         \add_1393/carry[15] , \add_1393/carry[14] , \add_1393/carry[13] ,
         \add_1393/carry[12] , \add_1393/carry[11] , \add_1393/carry[10] ,
         \add_1393/carry[9] , \add_1393/carry[8] , \add_1393/carry[7] ,
         \add_1393/carry[6] , \add_1393/carry[5] , \add_1393/carry[4] ,
         \add_1393/carry[3] , \add_1393/carry[2] , \add_1391/carry[31] ,
         \add_1391/carry[30] , \add_1391/carry[29] , \add_1391/carry[28] ,
         \add_1391/carry[27] , \add_1391/carry[26] , \add_1391/carry[25] ,
         \add_1391/carry[24] , \add_1391/carry[23] , \add_1391/carry[22] ,
         \add_1391/carry[21] , \add_1391/carry[20] , \add_1391/carry[19] ,
         \add_1391/carry[18] , \add_1391/carry[17] , \add_1391/carry[16] ,
         \add_1391/carry[15] , \add_1391/carry[14] , \add_1391/carry[13] ,
         \add_1391/carry[12] , \add_1391/carry[11] , \add_1391/carry[10] ,
         \add_1391/carry[9] , \add_1391/carry[8] , \add_1391/carry[7] ,
         \add_1391/carry[6] , \add_1391/carry[5] , \add_1391/carry[4] ,
         \add_1391/carry[3] , \add_1391/carry[2] , \add_1319/carry[31] ,
         \add_1319/carry[30] , \add_1319/carry[29] , \add_1319/carry[28] ,
         \add_1319/carry[27] , \add_1319/carry[26] , \add_1319/carry[25] ,
         \add_1319/carry[24] , \add_1319/carry[23] , \add_1319/carry[22] ,
         \add_1319/carry[21] , \add_1319/carry[20] , \add_1319/carry[19] ,
         \add_1319/carry[18] , \add_1319/carry[17] , \add_1319/carry[16] ,
         \add_1319/carry[15] , \add_1319/carry[14] , \add_1319/carry[13] ,
         \add_1319/carry[12] , \add_1319/carry[11] , \add_1319/carry[10] ,
         \add_1319/carry[9] , \add_1319/carry[8] , \add_1319/carry[7] ,
         \add_1319/carry[6] , \add_1319/carry[5] , \add_1319/carry[4] ,
         \add_1319/carry[3] , \add_1319/carry[2] , \sub_1275/carry[31] ,
         \sub_1275/carry[5] , \sub_1275/carry[4] , \sub_1275/carry[3] ,
         \sub_1275/carry[2] , \sub_1269/carry[31] , \sub_1269/carry[5] ,
         \sub_1269/carry[4] , \sub_1269/carry[3] , \sub_1269/carry[2] ,
         \sub_1263/carry[31] , \sub_1263/carry[5] , \sub_1263/carry[4] ,
         \sub_1263/carry[3] , \sub_1263/carry[2] , \sub_1255/carry[31] ,
         \sub_1255/carry[5] , \sub_1255/carry[4] , \sub_1255/carry[3] ,
         \sub_1255/carry[2] , \add_1125/carry[31] , \add_1125/carry[30] ,
         \add_1125/carry[29] , \add_1125/carry[28] , \add_1125/carry[27] ,
         \add_1125/carry[26] , \add_1125/carry[25] , \add_1125/carry[24] ,
         \add_1125/carry[23] , \add_1125/carry[22] , \add_1125/carry[21] ,
         \add_1125/carry[20] , \add_1125/carry[19] , \add_1125/carry[18] ,
         \add_1125/carry[17] , \add_1125/carry[16] , \add_1125/carry[15] ,
         \add_1125/carry[14] , \add_1125/carry[13] , \add_1125/carry[12] ,
         \add_1125/carry[11] , \add_1125/carry[10] , \add_1125/carry[9] ,
         \add_1125/carry[8] , \add_1125/carry[7] , \add_1125/carry[6] ,
         \add_1125/carry[5] , \add_1125/carry[4] , \add_1125/carry[3] ,
         \add_1125/carry[2] , \add_1121/carry[31] , \add_1121/carry[30] ,
         \add_1121/carry[29] , \add_1121/carry[28] , \add_1121/carry[27] ,
         \add_1121/carry[26] , \add_1121/carry[25] , \add_1121/carry[24] ,
         \add_1121/carry[23] , \add_1121/carry[22] , \add_1121/carry[21] ,
         \add_1121/carry[20] , \add_1121/carry[19] , \add_1121/carry[18] ,
         \add_1121/carry[17] , \add_1121/carry[16] , \add_1121/carry[15] ,
         \add_1121/carry[14] , \add_1121/carry[13] , \add_1121/carry[12] ,
         \add_1121/carry[11] , \add_1121/carry[10] , \add_1121/carry[9] ,
         \add_1121/carry[8] , \add_1121/carry[7] , \add_1121/carry[6] ,
         \add_1121/carry[5] , \add_1121/carry[4] , \add_1121/carry[3] ,
         \add_1121/carry[2] , n4688, n4689, n4690, n4691, n4692, n4693, n4694,
         n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704,
         n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724,
         n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734,
         n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744,
         n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754,
         n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764,
         n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774,
         n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784,
         n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794,
         n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804,
         n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814,
         n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824,
         n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834,
         n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874,
         n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884,
         n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894,
         n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904,
         n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914,
         n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924,
         n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934,
         n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944,
         n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954,
         n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964,
         n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974,
         n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984,
         n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994,
         n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004,
         n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014,
         n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024,
         n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034,
         n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044,
         n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054,
         n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084,
         n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094,
         n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104,
         n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114,
         n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124,
         n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134,
         n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144,
         n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154,
         n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164,
         n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174,
         n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184,
         n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194,
         n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204,
         n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214,
         n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224,
         n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234,
         n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244,
         n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254,
         n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264,
         n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274,
         n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284,
         n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294,
         n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304,
         n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314,
         n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344,
         n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354,
         n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364,
         n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374,
         n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384,
         n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394,
         n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404,
         n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414,
         n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424,
         n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434,
         n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444,
         n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454,
         n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464,
         n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474,
         n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484,
         n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494,
         n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504,
         n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514,
         n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524,
         n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554,
         n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564,
         n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574,
         n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584,
         n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594,
         n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604,
         n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614,
         n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624,
         n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634,
         n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644,
         n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654,
         n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664,
         n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674,
         n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684,
         n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694,
         n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704,
         n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714,
         n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724,
         n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734,
         n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744,
         n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754,
         n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764,
         n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774,
         n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784,
         n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794,
         n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804,
         n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814,
         n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824,
         n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834,
         n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844,
         n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854,
         n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864,
         n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874,
         n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884,
         n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894,
         n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904,
         n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914,
         n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924,
         n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934,
         n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944,
         n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954,
         n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964,
         n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974,
         n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984,
         n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994,
         n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004,
         n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014,
         n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024,
         n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034,
         n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044,
         n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054,
         n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064,
         n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074,
         n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084,
         n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094,
         n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104,
         n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114,
         n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124,
         n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134,
         n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144,
         n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154,
         n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164,
         n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174,
         n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184,
         n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194,
         n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204,
         n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214,
         n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224,
         n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234,
         n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264,
         n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274,
         n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284,
         n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294,
         n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304,
         n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314,
         n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324,
         n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354,
         n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364,
         n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374,
         n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384,
         n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394,
         n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404,
         n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414,
         n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424,
         n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434,
         n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444,
         n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454,
         n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464,
         n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474,
         n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484,
         n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494,
         n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504,
         n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514,
         n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524,
         n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534,
         n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544,
         n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554,
         n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564,
         n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574,
         n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584,
         n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594,
         n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604,
         n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614,
         n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674,
         n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684,
         n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694,
         n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704,
         n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714,
         n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724,
         n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734,
         n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744,
         n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754,
         n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764,
         n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774,
         n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784,
         n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794,
         n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804,
         n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814,
         n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824,
         n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834,
         n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844,
         n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854,
         n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864,
         n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874,
         n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884,
         n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894,
         n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904,
         n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914,
         n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924,
         n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934,
         n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964,
         n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974,
         n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984,
         n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994,
         n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004,
         n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014,
         n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024,
         n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034,
         n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044,
         n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054,
         n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064,
         n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074,
         n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084,
         n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094,
         n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104,
         n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114,
         n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124,
         n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134,
         n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144,
         n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194,
         n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204,
         n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214,
         n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224,
         n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234,
         n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244,
         n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254,
         n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264,
         n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274,
         n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284,
         n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294,
         n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304,
         n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314,
         n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324,
         n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334,
         n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344,
         n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354,
         n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364,
         n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374,
         n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384,
         n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394,
         n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404,
         n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444,
         n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454,
         n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464,
         n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474,
         n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484,
         n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494,
         n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504,
         n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514,
         n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524,
         n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534,
         n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564,
         n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574,
         n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584,
         n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594,
         n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604,
         n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614,
         n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644,
         n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654,
         n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664,
         n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674,
         n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684,
         n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694,
         n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704,
         n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714,
         n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724,
         n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734,
         n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744,
         n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754,
         n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764,
         n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774,
         n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784,
         n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794,
         n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804,
         n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814,
         n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824,
         n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834,
         n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844,
         n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854,
         n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864,
         n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874,
         n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884,
         n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894,
         n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904,
         n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914,
         n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944,
         n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954,
         n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964,
         n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974,
         n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984,
         n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994,
         n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004,
         n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014,
         n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024,
         n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034,
         n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044,
         n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054,
         n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064,
         n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074,
         n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084,
         n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094,
         n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104,
         n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114,
         n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124,
         n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134,
         n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144,
         n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154,
         n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164,
         n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174,
         n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184,
         n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194,
         n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204,
         n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214,
         n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224,
         n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234,
         n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244,
         n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254,
         n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264,
         n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274,
         n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284,
         n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294,
         n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304,
         n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314,
         n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324,
         n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334,
         n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344,
         n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354,
         n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364,
         n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374,
         n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384,
         n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394,
         n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404,
         n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414,
         n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424,
         n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434,
         n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444,
         n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454,
         n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464,
         n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474,
         n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484,
         n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494,
         n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504,
         n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514,
         n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524,
         n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534,
         n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544,
         n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554,
         n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564,
         n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574,
         n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584,
         n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594,
         n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604,
         n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614,
         n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624,
         n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634,
         n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644,
         n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654,
         n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664,
         n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674,
         n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684,
         n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694,
         n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704,
         n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714,
         n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724,
         n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734,
         n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744,
         n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754,
         n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764,
         n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774,
         n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784,
         n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794,
         n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804,
         n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814,
         n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824,
         n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834,
         n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844,
         n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854,
         n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864,
         n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874,
         n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884,
         n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894,
         n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904,
         n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914,
         n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924,
         n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934,
         n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944,
         n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954,
         n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964,
         n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974,
         n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984,
         n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994,
         n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004,
         n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014,
         n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024,
         n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034,
         n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044,
         n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054,
         n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064,
         n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074,
         n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084,
         n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094,
         n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104,
         n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114,
         n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124,
         n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134,
         n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144,
         n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154,
         n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164,
         n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174,
         n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184,
         n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194,
         n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204,
         n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214,
         n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224,
         n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234,
         n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244,
         n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254,
         n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264,
         n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274,
         n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284,
         n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294,
         n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304,
         n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314,
         n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324,
         n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334,
         n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344,
         n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354,
         n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364,
         n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374,
         n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384,
         n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394,
         n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404,
         n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414,
         n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424,
         n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434,
         n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444,
         n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454,
         n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464,
         n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474,
         n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484,
         n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494,
         n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504,
         n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514,
         n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524,
         n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534,
         n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544,
         n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554,
         n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564,
         n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574,
         n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584,
         n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594,
         n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604,
         n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614,
         n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624,
         n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634,
         n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644,
         n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654,
         n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664,
         n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674,
         n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684,
         n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694,
         n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704,
         n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714,
         n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724,
         n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734,
         n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744,
         n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754,
         n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764,
         n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774,
         n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784,
         n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794,
         n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804,
         n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814,
         n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824,
         n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834,
         n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844,
         n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854,
         n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864,
         n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874,
         n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884,
         n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894,
         n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904,
         n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914,
         n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924,
         n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934,
         n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944,
         n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954,
         n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964,
         n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974,
         n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984,
         n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994,
         n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003,
         n10004, n10005, n10006, n10007, n10008, n10009, n10010, n10011,
         n10012, n10013, n10014, n10015, n10016, n10017, n10018, n10019,
         n10020, n10021, n10022, n10023, n10024, n10025, n10026, n10027,
         n10028, n10029, n10030, n10031, n10032, n10033, n10034, n10035,
         n10036, n10037, n10038, n10039, n10040, n10041, n10042, n10043,
         n10044, n10045, n10046, n10047, n10048, n10049, n10050, n10051,
         n10052, n10053, n10054, n10055, n10056, n10057, n10058, n10059,
         n10060, n10061, n10062, n10063, n10064, n10065, n10066, n10067,
         n10068, n10069, n10070, n10071, n10072, n10073, n10074, n10075,
         n10076, n10077, n10078, n10079, n10080, n10081, n10082, n10083,
         n10084, n10085, n10086, n10087, n10088, n10089, n10090, n10091,
         n10092, n10093, n10094, n10095, n10096, n10097, n10098, n10099,
         n10100, n10101, n10102, n10103, n10104, n10105, n10106, n10107,
         n10108, n10109, n10110, n10111, n10112, n10113, n10114, n10115,
         n10116, n10117, n10118, n10119, n10120, n10121, n10122, n10123,
         n10124, n10125, n10126, n10127, n10128, n10129, n10130, n10131,
         n10132, n10133, n10134, n10135, n10136, n10137, n10138, n10139,
         n10140, n10141, n10142, n10143, n10144, n10145, n10146, n10147,
         n10148, n10149, n10150, n10151, n10152, n10153, n10154, n10155,
         n10156, n10157, n10158, n10159, n10160, n10161, n10162, n10163,
         n10164, n10165, n10166, n10167, n10168, n10169, n10170, n10171,
         n10172, n10173, n10174, n10175, n10176, n10177, n10178, n10179,
         n10180, n10181, n10182, n10183, n10184, n10185, n10186, n10187,
         n10188, n10189, n10190, n10191, n10192, n10193, n10194, n10195,
         n10196, n10197, n10198, n10199, n10200, n10201, n10202, n10203,
         n10204, n10205, n10206, n10207, n10208, n10209, n10210, n10211,
         n10212, n10213, n10214, n10215, n10216, n10217, n10218, n10219,
         n10220, n10221, n10222, n10223, n10224, n10225, n10226, n10227,
         n10228, n10229, n10230, n10231, n10232, n10233, n10234, n10235,
         n10236, n10237, n10238, n10239, n10240, n10241, n10242, n10243,
         n10244, n10245, n10246, n10247, n10248, n10249, n10250, n10251,
         n10252, n10253, n10254, n10255, n10256, n10257, n10258, n10259,
         n10260, n10261, n10262, n10263, n10264, n10265, n10266, n10267,
         n10268, n10269, n10270, n10271, n10272, n10273, n10274, n10275,
         n10276, n10277, n10278, n10279, n10280, n10281, n10282, n10283,
         n10284, n10285, n10286, n10287, n10288, n10289, n10290, n10291,
         n10292, n10293, n10294, n10295, n10296, n10297, n10298, n10299,
         n10300, n10301, n10302, n10303, n10304, n10305, n10306, n10307,
         n10308, n10309, n10310, n10311, n10312, n10313, n10314, n10315,
         n10316, n10317, n10318, n10319, n10320, n10321, n10322, n10323,
         n10324, n10325, n10326, n10327, n10328, n10329, n10330, n10331,
         n10332, n10333, n10334, n10335, n10336, n10337, n10338, n10339,
         n10340, n10341, n10342, n10343, n10344, n10345, n10346, n10347,
         n10348, n10349, n10350, n10351, n10352, n10353, n10354, n10355,
         n10356, n10357, n10358, n10359, n10360, n10361, n10362, n10363,
         n10364, n10365, n10366, n10367, n10368, n10369, n10370, n10371,
         n10372, n10373, n10374, n10375, n10376, n10377, n10378, n10379,
         n10380, n10381, n10382, n10383, n10384, n10385, n10386, n10387,
         n10388, n10389, n10390, n10391, n10392, n10393, n10394, n10395,
         n10396, n10397, n10398, n10399, n10400, n10401, n10402, n10403,
         n10404, n10405, n10406, n10407, n10408, n10409, n10410, n10411,
         n10412, n10413, n10414, n10415, n10416, n10417, n10418, n10419,
         n10420, n10421, n10422, n10423, n10424, n10425, n10426, n10427,
         n10428, n10429, n10430, n10431, n10432, n10433, n10434, n10435,
         n10436, n10437, n10438, n10439, n10440, n10441, n10442, n10443,
         n10444, n10445, n10446, n10447, n10448, n10449, n10450, n10451,
         n10452, n10453, n10454, n10455, n10456, n10457, n10458, n10459,
         n10460, n10461, n10462, n10463, n10464, n10465, n10466, n10467,
         n10468, n10469, n10470, n10471, n10472, n10473, n10474, n10475,
         n10476, n10477, n10478, n10479, n10480, n10481, n10482, n10483,
         n10484, n10485, n10486, n10487, n10488, n10489, n10490, n10491,
         n10492, n10493, n10494, n10495, n10496, n10497, n10498, n10499,
         n10500, n10501, n10502, n10503, n10504, n10505, n10506, n10507,
         n10508, n10509, n10510, n10511, n10512, n10513, n10514, n10515,
         n10516, n10517, n10518, n10519, n10520, n10521, n10522, n10523,
         n10524, n10525, n10526, n10527, n10528, n10529, n10530, n10531,
         n10532, n10533, n10534, n10535, n10536, n10537, n10538, n10539,
         n10540, n10541, n10542, n10543, n10544, n10545, n10546, n10547,
         n10548, n10549, n10550, n10551, n10552, n10553, n10554, n10555,
         n10556, n10557, n10558, n10559, n10560, n10561, n10562, n10563,
         n10564, n10565, n10566, n10567, n10568, n10569, n10570, n10571,
         n10572, n10573, n10574, n10575, n10576, n10577, n10578, n10579,
         n10580, n10581, n10582, n10583, n10584, n10585, n10586, n10587,
         n10588, n10589, n10590, n10591, n10592, n10593, n10594, n10595,
         n10596, n10597, n10598, n10599, n10600, n10601, n10602, n10603,
         n10604, n10605, n10606, n10607, n10608, n10609, n10610, n10611,
         n10612, n10613, n10614, n10615, n10616, n10617, n10618, n10619,
         n10620, n10621, n10622, n10623, n10624, n10625, n10626, n10627,
         n10628, n10629, n10630, n10631, n10632, n10633, n10634, n10635,
         n10636, n10637, n10638, n10639, n10640, n10641, n10642, n10643,
         n10644, n10645, n10646, n10647, n10648, n10649, n10650, n10651,
         n10652, n10653, n10654, n10655, n10656, n10657, n10658, n10659,
         n10660, n10661, n10662, n10663, n10664, n10665, n10666, n10667,
         n10668, n10669, n10670, n10671, n10672, n10673, n10674, n10675,
         n10676, n10677, n10678, n10679, n10680, n10681, n10682, n10683,
         n10684, n10685, n10686, n10687, n10688, n10689, n10690, n10691,
         n10692, n10693, n10694, n10695, n10696, n10697, n10698, n10699,
         n10700, n10701, n10702, n10703, n10704, n10705, n10706, n10707,
         n10708, n10709, n10710, n10711, n10712, n10713, n10714, n10715,
         n10716, n10717, n10718, n10719, n10720, n10721, n10722, n10723,
         n10724, n10725, n10726, n10727, n10728, n10729, n10730, n10731,
         n10732, n10733, n10734, n10735, n10736, n10737, n10738, n10739,
         n10740, n10741, n10742, n10743, n10744, n10745, n10746, n10747,
         n10748, n10749, n10750, n10751, n10752, n10753, n10754, n10755,
         n10756, n10757, n10758, n10759, n10760, n10761, n10762, n10763,
         n10764, n10765, n10766, n10767, n10768, n10769, n10770, n10771,
         n10772, n10773, n10774, n10775, n10776, n10777, n10778, n10779,
         n10780, n10781, n10782, n10783, n10784, n10785, n10786, n10787,
         n10788, n10789, n10790, n10791, n10792, n10793, n10794, n10795,
         n10796, n10797, n10798, n10799, n10800, n10801, n10802, n10803,
         n10804, n10805, n10806, n10807, n10808, n10809, n10810, n10811,
         n10812, n10813, n10814, n10815, n10816, n10817, n10818, n10819,
         n10820, n10821, n10822, n10823, n10824, n10825, n10826, n10827,
         n10828, n10829, n10830, n10831, n10832, n10833, n10834, n10835,
         n10836, n10837, n10838, n10839, n10840, n10841, n10842, n10843,
         n10844, n10845, n10846, n10847, n10848, n10849, n10850, n10851,
         n10852, n10853, n10854, n10855, n10856, n10857, n10858, n10859,
         n10860, n10861, n10862, n10863, n10864, n10865, n10866, n10867,
         n10868, n10869, n10870, n10871, n10872, n10873, n10874, n10875,
         n10876, n10877, n10878, n10879, n10880, n10881, n10882, n10883,
         n10884, n10885, n10886, n10887, n10888, n10889, n10890, n10892,
         n10893, n10894, n10895, n10896, n10897, n10898, n10899, n10900,
         n10901, n10902, n10903, n10904, n10905, n10906, n10907, n10908,
         n10909, n10910, n10911, n10912, n10913, n10914, n10915, n10916,
         n10917, n10918, n10919, n10920, n10921, n10922, n10923, n10924,
         n10925, n10926, n10927, n10928, n10929, n10930, n10931, n10932,
         n10933, n10934, n10935, n10936, n10937, n10938, n10939, n10940,
         n10941, n10942, n10943, n10944, n10945, n10946, n10947, n10948,
         n10949, n10950, n10951, n10952, n10953, n10954, n10955, n10956,
         n10957, n10958, n10959, n10960, n10961, n10962, n10963, n10964,
         n10965, n10966, n10967, n10968, n10969, n10970, n10971, n10972,
         n10973, n10974, n10975, n10976, n10977, n10978, n10979, n10980,
         n10981, n10982, n10983, n10984, n10985, n10986, n10987, n10988,
         n10989, n10990, n10991, n10992, n10993, n10994, n10995, n10996,
         n10997, n10998, n10999, n11000, n11001, n11002, n11003, n11004,
         n11005, n11006, n11007, n11008, n11009, n11010, n11011, n11012,
         n11013, n11014, n11015, n11016, n11017, n11018, n11019, n11020,
         n11021, n11022, n11023, n11024, n11025, n11026, n11027, n11028,
         n11029, n11030, n11031, n11032, n11033, n11034, n11035, n11036,
         n11037, n11038, n11039, n11040, n11041, n11042, n11043, n11044,
         n11045, n11046, n11047, n11048, n11049, n11050, n11051, n11052,
         n11053, n11054, n11055, n11056, n11057, n11058, n11059, n11060,
         n11061, n11062, n11063, n11064, n11065, n11066, n11067, n11068,
         n11069, n11070, n11071, n11072, n11073, n11074, n11075, n11076,
         n11077, n11078, n11079, n11080, n11081, n11082, n11083, n11084,
         n11085, n11086, n11087, n11088, n11089, n11090, n11091, n11092,
         n11093, n11094, n11095, n11096, n11097, n11098, n11099, n11100,
         n11101, n11102, n11103, n11104, n11105, n11106, n11107, n11108,
         n11109, n11110, n11111, n11112, n11113, n11114, n11115, n11116,
         n11117, n11118, n11119, n11120, n11121, n11122, n11123, n11124,
         n11125, n11126, n11127, n11128, n11129, n11130, n11131, n11132,
         n11133, n11134, n11135, n11136, n11137, n11138, n11139, n11140,
         n11141, n11142, n11143, n11144, n11145, n11146, n11147, n11148,
         n11149, n11150, n11151, n11152, n11153, n11154, n11155, n11156,
         n11157, n11158, n11159, n11160, n11161, n11162, n11163, n11164,
         n11165, n11166, n11167, n11168, n11169, n11170, n11171, n11172,
         n11173, n11174, n11175, n11176, n11177, n11178, n11179, n11180,
         n11181, n11182, n11183, n11184, n11185, n11186, n11187, n11188,
         n11189, n11190, n11191, n11192, n11193, n11194, n11195, n11196,
         n11197, n11198, n11199, n11200, n11201, n11202, n11203, n11204,
         n11205, n11206, n11207, n11208, n11209, n11210, n11211, n11212,
         n11213, n11214, n11215, n11216, n11217, n11218, n11219, n11220,
         n11221, n11222, n11223, n11224, n11225, n11226, n11227, n11228,
         n11229, n11230, n11231, n11232, n11233, n11234, n11235, n11236,
         n11237, n11238, n11239, n11240, n11241, n11242, n11243, n11244,
         n11245, n11246, n11247, n11248, n11249, n11250, n11251, n11252,
         n11253, n11254, n11255, n11256, n11257, n11258, n11259, n11260,
         n11261, n11262, n11263, n11264, n11265, n11266, n11267, n11268,
         n11269, n11270, n11271, n11272, n11273, n11274, n11275, n11276,
         n11277, n11278, n11279, n11280, n11281, n11282, n11283, n11284,
         n11285, n11286, n11287, n11288, n11289, n11290, n11291, n11292,
         n11293, n11294, n11295, n11296, n11297, n11298, n11299, n11300,
         n11301, n11302, n11303, n11304, n11305, n11306, n11307, n11308,
         n11309, n11310, n11311, n11312, n11313, n11314, n11315, n11316,
         n11317, n11318, n11319, n11320, n11321, n11322, n11323, n11324,
         n11325, n11326, n11327, n11328, n11329, n11330, n11331, n11332,
         n11333, n11334, n11335, n11336, n11337, n11338, n11339, n11340,
         n11341, n11342, n11343, n11344, n11345, n11346, n11347, n11348,
         n11349, n11350, n11351, n11352, n11353, n11354, n11355, n11356,
         n11357, n11358, n11359, n11360, n11361, n11362, n11363, n11364,
         n11365, n11366, n11367, n11368, n11369, n11370, n11371, n11372,
         n11373, n11374, n11375, n11376, n11377, n11378, n11379, n11380,
         n11381, n11382, n11383, n11384, n11385, n11386, n11387, n11388,
         n11389, n11390, n11391, n11392, n11393, n11394, n11395, n11396,
         n11397, n11398, n11399, n11400, n11401, n11402, n11403, n11404,
         n11405, n11406, n11407, n11408, n11409, n11410, n11411, n11412,
         n11413, n11414, n11415, n11416, n11417, n11418, n11419, n11420,
         n11421, n11422, n11423, n11424, n11425, n11426, n11427, n11428,
         n11429, n11430, n11431, n11432, n11433, n11434, n11435, n11436,
         n11437, n11438, n11439, n11440, n11441, n11442, n11443, n11444,
         n11445, n11446, n11447, n11448, n11449, n11450, n11451, n11452,
         n11453, n11454, n11455, n11456, n11457, n11458, n11459, n11460,
         n11461, n11462, n11463, n11464, n11465, n11466, n11467, n11468,
         n11469, n11470, n11471, n11472, n11473, n11474, n11475, n11476,
         n11477, n11478, n11479, n11480, n11481, n11482, n11483, n11484,
         n11485, n11486, n11487, n11488, n11489, n11490, n11491, n11492,
         n11493, n11494, n11495, n11496, n11497, n11498, n11499, n11500,
         n11501, n11502, n11503, n11504, n11505, n11506, n11507, n11508,
         n11509, n11510, n11511, n11512, n11513, n11514, n11515, n11516,
         n11517, n11518, n11519, n11520, n11521, n11522, n11523, n11524,
         n11525, n11526, n11527, n11528, n11529, n11530, n11531, n11532,
         n11533, n11534, n11535, n11536, n11537, n11538, n11539, n11540,
         n11541, n11542, n11543, n11544, n11545, n11546, n11547, n11548,
         n11549, n11550, n11551, n11552, n11553, n11554, n11555, n11556,
         n11557, n11558, n11559, n11560, n11561, n11562, n11563, n11564,
         n11565, n11566, n11567, n11568, n11569, n11570, n11571, n11572,
         n11573, n11574, n11575, n11576, n11577, n11578, n11579, n11580,
         n11581, n11582, n11583, n11584, n11585, n11586, n11587, n11588,
         n11589, n11590, n11591, n11592, n11593, n11594, n11595, n11596,
         n11597, n11598, n11599, n11600, n11601, n11602, n11603, n11604,
         n11605, n11606, n11607, n11608, n11609, n11610, n11611, n11612,
         n11613, n11614, n11615, n11616, n11617, n11618, n11619, n11620,
         n11621, n11622, n11623, n11624, n11625, n11626, n11627, n11628,
         n11629, n11630, n11631, n11632, n11633, n11634, n11635, n11636,
         n11637, n11638, n11639, n11640, n11641, n11642, n11643, n11644,
         n11645, n11646, n11647, n11648, n11649, n11650, n11651, n11652,
         n11653, n11654, n11655, n11656, n11657, n11658, n11659, n11660,
         n11661, n11662, n11663, n11664, n11665, n11666, n11667, n11668,
         n11669, n11670, n11671, n11672, n11673, n11674, n11675, n11676,
         n11677, n11678, n11679, n11680, n11681, n11682, n11683, n11684,
         n11685, n11686, n11687, n11688, n11689, n11690, n11691, n11692,
         n11693, n11694, n11695, n11696, n11697, n11698, n11699, n11700,
         n11701, n11702, n11703, n11704, n11705, n11706, n11707, n11708,
         n11709, n11710, n11711, n11712, n11713, n11714, n11715, n11716,
         n11717, n11718, n11719, n11720, n11721, n11722, n11723, n11724,
         n11725, n11726, n11727, n11728, n11729, n11730, n11731, n11732,
         n11733, n11734, n11735, n11736, n11737, n11738, n11739, n11740,
         n11741, n11742, n11743, n11744, n11745, n11746, n11747, n11748,
         n11749, n11750, n11751, n11752, n11753, n11754, n11755, n11756,
         n11757, n11758, n11759, n11760, n11761, n11762, n11763, n11764,
         n11765, n11766, n11767, n11768, n11769, n11770, n11771, n11772,
         n11773, n11774, n11775, n11776, n11777, n11778, n11779, n11780,
         n11781, n11782, n11783, n11784, n11785, n11786, n11787, n11788,
         n11789, n11790, n11791, n11792, n11793, n11794, n11795, n11796,
         n11797, n11798, n11799, n11800, n11801, n11802, n11803, n11804,
         n11805, n11806, n11807, n11808, n11809, n11810, n11811, n11812,
         n11813, n11814, n11815, n11816, n11817, n11818, n11819, n11820,
         n11821, n11822, n11823, n11824, n11825, n11826, n11827, n11828,
         n11829, n11830, n11831, n11832, n11833, n11834, n11835, n11836,
         n11837, n11838, n11839, n11840, n11841, n11842, n11843, n11844,
         n11845, n11846, n11847, n11848, n11849, n11850, n11851, n11852,
         n11853, n11854, n11855, n11856, n11857, n11858, n11859, n11860,
         n11861, n11862, n11863, n11864, n11865, n11866, n11867, n11868,
         n11869, n11870, n11871, n11872, n11873, n11874, n11875, n11876,
         n11877, n11878, n11879, n11880, n11881, n11882, n11883, n11884,
         n11885, n11886, n11887, n11888, n11889, n11890, n11891, n11892,
         n11893, n11894, n11895, n11896, n11897, n11898, n11899, n11900,
         n11901, n11902, n11903, n11904, n11905, n11906, n11907, n11908,
         n11909, n11910, n11911, n11912, n11913, n11914, n11915, n11916,
         n11917, n11918, n11919, n11920, n11921, n11922, n11923, n11924,
         n11925, n11926, n11927, n11928, n11929, n11930, n11931, n11932,
         n11933, n11934, n11935, n11936, n11937, n11938, n11939, n11940,
         n11941, n11942, n11943, n11944, n11945, n11946, n11947, n11948,
         n11949, n11950, n11951, n11952, n11953, n11954, n11955, n11956,
         n11957, n11958, n11959, n11960, n11961, n11962, n11963, n11964,
         n11965, n11966, n11967, n11968, n11969, n11970, n11971, n11972,
         n11973, n11974, n11975, n11976, n11977, n11978, n11979, n11980,
         n11981, n11982, n11983, n11984, n11985, n11986, n11987, n11988,
         n11989, n11990, n11991, n11992, n11993, n11994, n11995, n11996,
         n11997, n11998, n11999, n12000, n12001, n12002, n12003, n12004,
         n12005, n12006, n12007, n12008, n12009, n12010, n12011, n12012,
         n12013, n12014, n12015, n12016, n12017, n12018, n12019, n12020,
         n12021, n12022, n12023, n12024, n12025, n12026, n12027, n12028,
         n12029, n12030, n12031, n12032, n12033, n12034, n12035, n12036,
         n12037, n12038, n12039, n12040, n12041, n12042, n12043, n12044,
         n12045, n12046, n12047, n12048, n12049, n12050, n12051, n12052,
         n12053, n12054, n12055, n12056, n12057, n12058, n12059, n12060,
         n12061, n12062, n12063, n12064, n12065, n12066, n12067, n12068,
         n12069, n12070, n12071, n12072, n12073, n12074, n12075, n12076,
         n12077, n12078, n12079, n12080, n12081, n12082, n12083, n12084,
         n12085, n12086, n12087, n12088, n12089, n12090, n12091, n12092,
         n12093, n12094, n12095, n12096, n12097, n12098, n12099, n12100,
         n12101, n12102, n12103, n12104, n12105, n12106, n12107, n12108,
         n12109, n12110, n12111, n12112, n12113, n12114, n12115, n12116,
         n12117, n12118, n12119, n12120, n12121, n12122, n12123, n12124,
         n12125, n12126, n12127, n12128, n12129, n12130, n12131, n12132,
         n12133, n12134, n12135, n12136, n12137, n12138, n12139, n12140,
         n12141, n12142, n12143, n12144, n12145, n12146, n12147, n12148,
         n12149, n12150, n12151, n12152, n12153, n12154, n12155, n12156,
         n12157, n12158, n12159, n12160, n12161, n12162, n12163, n12164,
         n12165, n12166, n12167, n12168, n12169, n12170, n12171, n12172,
         n12173, n12174, n12175, n12176, n12177, n12178, n12179, n12180,
         n12181, n12182, n12183, n12184, n12185, n12186, n12187, n12188,
         n12189, n12190, n12191, n12192, n12193, n12194, n12195, n12196,
         n12197, n12198, n12199, n12200, n12201, n12202, n12203, n12204,
         n12205, n12206, n12207, n12208, n12209, n12210, n12211, n12212,
         n12213, n12214, n12215, n12216, n12217, n12218, n12219, n12220,
         n12221, n12222, n12223, n12224, n12225, n12226, n12227, n12228,
         n12229, n12230, n12231, n12232, n12233, n12234, n12235, n12236,
         n12237, n12238, n12239, n12240, n12241, n12242, n12243, n12244,
         n12245, n12246, n12247, n12248, n12249, n12250, n12251, n12252,
         n12253, n12254, n12255, n12256, n12257, n12258, n12259, n12260,
         n12261, n12262, n12263, n12264;
  wire   [4:0] recentdatapoints_data_address0;
  wire   [15:0] data_read_reg_1495;
  wire   [15:0] recentdatapoints_data_q0;
  wire   [4:0] recentVBools_data_address0;
  wire   [4:0] recentABools_data_address0;
  wire   [31:0] athresh;
  wire   [31:0] vthresh;
  wire   [7:0] a_flip;
  wire   [7:0] v_flip;
  wire   [31:0] a_length;
  wire   [31:0] v_length;
  wire   [15:0] data;
  wire   [13:0] ap_CS_fsm;
  wire   [31:0] ACaptureThresh_loc_reg_288;
  wire   [31:0] ACaptureThresh;
  wire   [31:0] AbeatDelay_new_reg_394;
  wire   [31:0] tmp_3_reg_1589;
  wire   [31:0] VCaptureThresh_loc_reg_298;
  wire   [31:0] VCaptureThresh;
  wire   [31:0] VbeatDelay_new_1_reg_326;
  wire   [31:0] tmp_4_reg_1596;
  wire   [31:0] VbeatFallDelay_new_1_reg_342;
  wire   [31:0] tmp_5_reg_1603;
  wire   [31:0] recentABools_len_new_reg_385;
  wire   [31:0] CircularBuffer_len_read_assign_3_fu_1091_p3;
  wire   [31:0] CircularBuffer_len_write_assig_3_fu_1249_p2;
  wire   [31:0] recentVBools_len_new_reg_317;
  wire   [31:0] CircularBuffer_len_read_assign_1_fu_778_p3;
  wire   [31:0] CircularBuffer_len_write_assig_1_fu_924_p2;
  wire   [31:0] sum_1_reg_376;
  wire   [31:0] CircularBuffer_sum_write_assig_3_fu_1242_p2;
  wire   [31:0] sum_reg_308;
  wire   [31:0] CircularBuffer_sum_write_assig_1_fu_917_p2;
  wire   [31:0] a_thresh;
  wire   [7:0] aflip;
  wire   [31:0] v_thresh;
  wire   [7:0] vflip;
  wire   [31:0] AbeatDelay;
  wire   [31:0] AstimDelay;
  wire   [31:0] VstimDelay;
  wire   [31:0] CircularBuffer_head_i_read_ass_1_fu_1110_p3;
  wire   [31:0] CircularBuffer_head_i_read_ass_1_reg_1719;
  wire   [31:0] CircularBuffer_len_read_assign_3_reg_1711;
  wire   [31:0] CircularBuffer_sum_read_assign_1_reg_1705;
  wire   [31:0] VbeatDelay;
  wire   [31:0] VbeatFallDelay;
  wire   [31:0] recentABools_head_i;
  wire   [31:0] CircularBuffer_head_i_read_ass_fu_797_p3;
  wire   [31:0] CircularBuffer_head_i_read_ass_reg_1624;
  wire   [31:0] CircularBuffer_len_read_assign_1_reg_1616;
  wire   [31:0] CircularBuffer_sum_read_assign_reg_1610;
  wire   [31:0] recentVBools_head_i;
  wire   [31:0] tmp_3_fu_706_p2;
  wire   [31:0] tmp_4_fu_716_p2;
  wire   [31:0] tmp_5_fu_726_p2;
  wire   [31:0] CircularBuffer_len_write_assig_2_reg_1729;
  wire   [31:0] CircularBuffer_len_write_assig_2_fu_1142_p2;
  wire   [31:0] CircularBuffer_len_write_assig_reg_1634;
  wire   [31:0] CircularBuffer_len_write_assig_fu_817_p2;
  wire   [4:0] recentdatapoints_data_addr_reg_1533;
  wire   [31:0] tmp_6_reg_1538;
  wire   [31:0] tmp_6_fu_497_p3;
  wire   [31:0] tmp_7_reg_1544;
  wire   [31:0] tmp_7_fu_511_p3;
  wire   [31:0] p_tmp_i_fu_587_p3;
  wire   [31:0] p_tmp_i_reg_1556;
  wire   [31:0] recentdatapoints_head_i;
  wire   [31:0] recentdatapoints_len;
  wire   [31:0] tmp_38_i_reg_1550;
  wire   [4:0] recentABools_data_addr_reg_1689;
  wire   [31:0] recentVBools_len;
  wire   [31:0] recentVBools_sum;
  wire   [31:0] sum_phi_fu_311_p4;
  wire   [31:0] recentABools_len;
  wire   [31:0] recentABools_sum;
  wire   [31:0] sum_1_phi_fu_379_p4;
  wire   [4:0] recentVBools_data_addr_reg_1573;
  wire   [31:0] tmp_33_i1_fu_1099_p2;
  wire   [31:0] tmp_33_i_fu_786_p2;
  wire   [31:0] CircularBuffer_int_30_sum_i1_fu_1071_p3;
  wire   [31:0] tmp_29_i1_fu_1065_p2;
  wire   [31:0] CircularBuffer_int_30_sum_i_fu_758_p3;
  wire   [31:0] tmp_29_i_fu_752_p2;
  wire   [31:0] CircularBuffer_len_read_assign_fu_772_p2;
  wire   [31:0] CircularBuffer_len_read_assign_2_fu_1085_p2;
  wire   [16:0] datapointA_1_fu_1017_p2;
  wire   [16:0] datapointV_1_fu_674_p2;
  wire   [4:0] i_9_fu_1160_p2;
  wire   [31:0] i_8_fu_1148_p2;
  wire   [31:0] i_11_fu_1179_p2;
  wire   [4:0] i_12_fu_1191_p2;
  wire   [4:0] i_1_fu_620_p2;
  wire   [31:0] i_2_fu_823_p2;
  wire   [4:0] i_3_fu_835_p2;
  wire   [31:0] i_5_fu_854_p2;
  wire   [4:0] i_6_fu_866_p2;
  wire   [4:0] i_fu_607_p2;
  wire   [15:0] p_1_cast_fu_1031_p1;
  wire   [15:0] p_cast_fu_688_p1;
  wire   [31:0] tmp_39_i_fu_576_p2;
  wire   [31:0] recentdatapoints_len_load_op_fu_556_p2;
  assign s_axi_AXILiteS_RVALID = \Decision_AXILiteS_s_axi_U/rstate[0] ;
  assign s_axi_AXILiteS_BRESP[1] = 1'b0;
  assign s_axi_AXILiteS_BRESP[0] = 1'b0;
  assign s_axi_AXILiteS_RRESP[1] = 1'b0;
  assign s_axi_AXILiteS_RRESP[0] = 1'b0;

  DFFPOSX1 \toReturn_8_reg_1755_reg[0]  ( .D(n8218), .CLK(n9222), .Q(
        \toReturn_8_reg_1755[0] ) );
  DFFPOSX1 \recentABools_sum_reg[31]  ( .D(n4373), .CLK(n9222), .Q(
        recentABools_sum[31]) );
  DFFPOSX1 \sum_1_reg_376_reg[30]  ( .D(n4278), .CLK(n9222), .Q(
        sum_1_reg_376[30]) );
  DFFPOSX1 \tmp_19_reg_409_reg[0]  ( .D(n4168), .CLK(n9222), .Q(
        \tmp_19_reg_409[0] ) );
  DFFPOSX1 \ap_CS_fsm_reg[0]  ( .D(n4761), .CLK(n9222), .Q(ap_CS_fsm[0]) );
  DFFPOSX1 \aflip_reg[3]  ( .D(n4679), .CLK(n9222), .Q(aflip[3]) );
  DFFPOSX1 \aflip_reg[4]  ( .D(n4678), .CLK(n9221), .Q(aflip[4]) );
  DFFPOSX1 \aflip_reg[5]  ( .D(n4677), .CLK(n9221), .Q(aflip[5]) );
  DFFPOSX1 \aflip_reg[6]  ( .D(n4676), .CLK(n9221), .Q(aflip[6]) );
  DFFPOSX1 \aflip_reg[7]  ( .D(n4675), .CLK(n9221), .Q(aflip[7]) );
  DFFPOSX1 \v_thresh_reg[0]  ( .D(n9402), .CLK(n9221), .Q(v_thresh[0]) );
  DFFPOSX1 \v_thresh_reg[1]  ( .D(n9403), .CLK(n9221), .Q(v_thresh[1]) );
  DFFPOSX1 \v_thresh_reg[2]  ( .D(n9404), .CLK(n9221), .Q(v_thresh[2]) );
  DFFPOSX1 \v_thresh_reg[3]  ( .D(n9405), .CLK(n9221), .Q(v_thresh[3]) );
  DFFPOSX1 \v_thresh_reg[4]  ( .D(n9406), .CLK(n9221), .Q(v_thresh[4]) );
  DFFPOSX1 \v_thresh_reg[5]  ( .D(n9407), .CLK(n9221), .Q(v_thresh[5]) );
  DFFPOSX1 \v_thresh_reg[6]  ( .D(n9408), .CLK(n9221), .Q(v_thresh[6]) );
  DFFPOSX1 \v_thresh_reg[7]  ( .D(n9409), .CLK(n9221), .Q(v_thresh[7]) );
  DFFPOSX1 \v_thresh_reg[8]  ( .D(n9410), .CLK(n9221), .Q(v_thresh[8]) );
  DFFPOSX1 \v_thresh_reg[9]  ( .D(n9411), .CLK(n9220), .Q(v_thresh[9]) );
  DFFPOSX1 \v_thresh_reg[10]  ( .D(n9412), .CLK(n9220), .Q(v_thresh[10]) );
  DFFPOSX1 \v_thresh_reg[11]  ( .D(n9413), .CLK(n9220), .Q(v_thresh[11]) );
  DFFPOSX1 \v_thresh_reg[12]  ( .D(n9414), .CLK(n9220), .Q(v_thresh[12]) );
  DFFPOSX1 \v_thresh_reg[13]  ( .D(n9415), .CLK(n9220), .Q(v_thresh[13]) );
  DFFPOSX1 \v_thresh_reg[14]  ( .D(n9416), .CLK(n9220), .Q(v_thresh[14]) );
  DFFPOSX1 \v_thresh_reg[15]  ( .D(n9417), .CLK(n9220), .Q(v_thresh[15]) );
  DFFPOSX1 \v_thresh_reg[16]  ( .D(n9418), .CLK(n9220), .Q(v_thresh[16]) );
  DFFPOSX1 \v_thresh_reg[17]  ( .D(n9419), .CLK(n9220), .Q(v_thresh[17]) );
  DFFPOSX1 \v_thresh_reg[18]  ( .D(n9420), .CLK(n9220), .Q(v_thresh[18]) );
  DFFPOSX1 \v_thresh_reg[19]  ( .D(n9421), .CLK(n9220), .Q(v_thresh[19]) );
  DFFPOSX1 \v_thresh_reg[20]  ( .D(n9422), .CLK(n9220), .Q(v_thresh[20]) );
  DFFPOSX1 \v_thresh_reg[21]  ( .D(n9423), .CLK(n9220), .Q(v_thresh[21]) );
  DFFPOSX1 \v_thresh_reg[22]  ( .D(n9424), .CLK(n9219), .Q(v_thresh[22]) );
  DFFPOSX1 \v_thresh_reg[23]  ( .D(n9425), .CLK(n9219), .Q(v_thresh[23]) );
  DFFPOSX1 \v_thresh_reg[24]  ( .D(n9426), .CLK(n9219), .Q(v_thresh[24]) );
  DFFPOSX1 \v_thresh_reg[25]  ( .D(n9427), .CLK(n9219), .Q(v_thresh[25]) );
  DFFPOSX1 \v_thresh_reg[26]  ( .D(n9428), .CLK(n9219), .Q(v_thresh[26]) );
  DFFPOSX1 \v_thresh_reg[27]  ( .D(n9429), .CLK(n9219), .Q(v_thresh[27]) );
  DFFPOSX1 \v_thresh_reg[28]  ( .D(n9430), .CLK(n9219), .Q(v_thresh[28]) );
  DFFPOSX1 \v_thresh_reg[29]  ( .D(n9431), .CLK(n9219), .Q(v_thresh[29]) );
  DFFPOSX1 \v_thresh_reg[30]  ( .D(n9432), .CLK(n9219), .Q(v_thresh[30]) );
  DFFPOSX1 \v_thresh_reg[31]  ( .D(n9433), .CLK(n9219), .Q(v_thresh[31]) );
  DFFPOSX1 \vflip_reg[0]  ( .D(n4674), .CLK(n9219), .Q(vflip[0]) );
  DFFPOSX1 \vflip_reg[1]  ( .D(n4673), .CLK(n9219), .Q(vflip[1]) );
  DFFPOSX1 \vflip_reg[2]  ( .D(n4672), .CLK(n9219), .Q(vflip[2]) );
  DFFPOSX1 \vflip_reg[3]  ( .D(n4671), .CLK(n9218), .Q(vflip[3]) );
  DFFPOSX1 \vflip_reg[4]  ( .D(n4670), .CLK(n9218), .Q(vflip[4]) );
  DFFPOSX1 \vflip_reg[5]  ( .D(n4669), .CLK(n9218), .Q(vflip[5]) );
  DFFPOSX1 \vflip_reg[6]  ( .D(n4668), .CLK(n9218), .Q(vflip[6]) );
  DFFPOSX1 \vflip_reg[7]  ( .D(n4667), .CLK(n9218), .Q(vflip[7]) );
  DFFPOSX1 \ACaptureThresh_reg[0]  ( .D(n4666), .CLK(n9218), .Q(
        ACaptureThresh[0]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[0]  ( .D(n4771), .CLK(n9218), .Q(
        ACaptureThresh_loc_reg_288[0]) );
  DFFPOSX1 \ACaptureThresh_reg[1]  ( .D(n4665), .CLK(n9218), .Q(
        ACaptureThresh[1]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[1]  ( .D(n4772), .CLK(n9218), .Q(
        ACaptureThresh_loc_reg_288[1]) );
  DFFPOSX1 \ACaptureThresh_reg[2]  ( .D(n4664), .CLK(n9218), .Q(
        ACaptureThresh[2]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[2]  ( .D(n4773), .CLK(n9218), .Q(
        ACaptureThresh_loc_reg_288[2]) );
  DFFPOSX1 \ACaptureThresh_reg[3]  ( .D(n4663), .CLK(n9218), .Q(
        ACaptureThresh[3]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[3]  ( .D(n6086), .CLK(n9218), .Q(
        ACaptureThresh_loc_reg_288[3]) );
  DFFPOSX1 \ACaptureThresh_reg[4]  ( .D(n4662), .CLK(n9217), .Q(
        ACaptureThresh[4]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[4]  ( .D(n6240), .CLK(n9217), .Q(
        ACaptureThresh_loc_reg_288[4]) );
  DFFPOSX1 \ACaptureThresh_reg[5]  ( .D(n4661), .CLK(n9217), .Q(
        ACaptureThresh[5]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[5]  ( .D(n6335), .CLK(n9217), .Q(
        ACaptureThresh_loc_reg_288[5]) );
  DFFPOSX1 \ACaptureThresh_reg[6]  ( .D(n4660), .CLK(n9217), .Q(
        ACaptureThresh[6]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[6]  ( .D(n6444), .CLK(n9217), .Q(
        ACaptureThresh_loc_reg_288[6]) );
  DFFPOSX1 \ACaptureThresh_reg[7]  ( .D(n4659), .CLK(n9217), .Q(
        ACaptureThresh[7]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[7]  ( .D(n6557), .CLK(n9217), .Q(
        ACaptureThresh_loc_reg_288[7]) );
  DFFPOSX1 \ACaptureThresh_reg[8]  ( .D(n4658), .CLK(n9217), .Q(
        ACaptureThresh[8]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[8]  ( .D(n6666), .CLK(n9217), .Q(
        ACaptureThresh_loc_reg_288[8]) );
  DFFPOSX1 \ACaptureThresh_reg[9]  ( .D(n4657), .CLK(n9217), .Q(
        ACaptureThresh[9]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[9]  ( .D(n6155), .CLK(n9217), .Q(
        ACaptureThresh_loc_reg_288[9]) );
  DFFPOSX1 \ACaptureThresh_reg[10]  ( .D(n4656), .CLK(n9217), .Q(
        ACaptureThresh[10]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[10]  ( .D(n6787), .CLK(n9216), .Q(
        ACaptureThresh_loc_reg_288[10]) );
  DFFPOSX1 \ACaptureThresh_reg[11]  ( .D(n4655), .CLK(n9216), .Q(
        ACaptureThresh[11]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[11]  ( .D(n6922), .CLK(n9216), .Q(
        ACaptureThresh_loc_reg_288[11]) );
  DFFPOSX1 \ACaptureThresh_reg[12]  ( .D(n4654), .CLK(n9216), .Q(
        ACaptureThresh[12]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[12]  ( .D(n7983), .CLK(n9216), .Q(
        ACaptureThresh_loc_reg_288[12]) );
  DFFPOSX1 \ACaptureThresh_reg[13]  ( .D(n4653), .CLK(n9216), .Q(
        ACaptureThresh[13]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[13]  ( .D(n7065), .CLK(n9216), .Q(
        ACaptureThresh_loc_reg_288[13]) );
  DFFPOSX1 \ACaptureThresh_reg[14]  ( .D(n4652), .CLK(n9216), .Q(
        ACaptureThresh[14]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[14]  ( .D(n7221), .CLK(n9216), .Q(
        ACaptureThresh_loc_reg_288[14]) );
  DFFPOSX1 \ACaptureThresh_reg[15]  ( .D(n4651), .CLK(n9216), .Q(
        ACaptureThresh[15]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[15]  ( .D(n7386), .CLK(n9216), .Q(
        ACaptureThresh_loc_reg_288[15]) );
  DFFPOSX1 \ACaptureThresh_reg[16]  ( .D(n4650), .CLK(n9216), .Q(
        ACaptureThresh[16]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[16]  ( .D(n7571), .CLK(n9216), .Q(
        ACaptureThresh_loc_reg_288[16]) );
  DFFPOSX1 \ACaptureThresh_reg[17]  ( .D(n4649), .CLK(n9215), .Q(
        ACaptureThresh[17]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[17]  ( .D(n7765), .CLK(n9215), .Q(
        ACaptureThresh_loc_reg_288[17]) );
  DFFPOSX1 \ACaptureThresh_reg[18]  ( .D(n4648), .CLK(n9215), .Q(
        ACaptureThresh[18]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[18]  ( .D(n8224), .CLK(n9215), .Q(
        ACaptureThresh_loc_reg_288[18]) );
  DFFPOSX1 \ACaptureThresh_reg[19]  ( .D(n4647), .CLK(n9215), .Q(
        ACaptureThresh[19]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[19]  ( .D(n6158), .CLK(n9215), .Q(
        ACaptureThresh_loc_reg_288[19]) );
  DFFPOSX1 \ACaptureThresh_reg[20]  ( .D(n4646), .CLK(n9215), .Q(
        ACaptureThresh[20]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[20]  ( .D(n6243), .CLK(n9215), .Q(
        ACaptureThresh_loc_reg_288[20]) );
  DFFPOSX1 \ACaptureThresh_reg[21]  ( .D(n4645), .CLK(n9215), .Q(
        ACaptureThresh[21]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[21]  ( .D(n6338), .CLK(n9215), .Q(
        ACaptureThresh_loc_reg_288[21]) );
  DFFPOSX1 \ACaptureThresh_reg[22]  ( .D(n4644), .CLK(n9215), .Q(
        ACaptureThresh[22]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[22]  ( .D(n6447), .CLK(n9215), .Q(
        ACaptureThresh_loc_reg_288[22]) );
  DFFPOSX1 \ACaptureThresh_reg[23]  ( .D(n4643), .CLK(n9215), .Q(
        ACaptureThresh[23]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[23]  ( .D(n6560), .CLK(n9214), .Q(
        ACaptureThresh_loc_reg_288[23]) );
  DFFPOSX1 \ACaptureThresh_reg[24]  ( .D(n4642), .CLK(n9214), .Q(
        ACaptureThresh[24]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[24]  ( .D(n6669), .CLK(n9214), .Q(
        ACaptureThresh_loc_reg_288[24]) );
  DFFPOSX1 \ACaptureThresh_reg[25]  ( .D(n4641), .CLK(n9214), .Q(
        ACaptureThresh[25]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[25]  ( .D(n7986), .CLK(n9214), .Q(
        ACaptureThresh_loc_reg_288[25]) );
  DFFPOSX1 \ACaptureThresh_reg[26]  ( .D(n4640), .CLK(n9214), .Q(
        ACaptureThresh[26]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[26]  ( .D(n6790), .CLK(n9214), .Q(
        ACaptureThresh_loc_reg_288[26]) );
  DFFPOSX1 \ACaptureThresh_reg[27]  ( .D(n4639), .CLK(n9214), .Q(
        ACaptureThresh[27]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[27]  ( .D(n6925), .CLK(n9214), .Q(
        ACaptureThresh_loc_reg_288[27]) );
  DFFPOSX1 \ACaptureThresh_reg[28]  ( .D(n4638), .CLK(n9214), .Q(
        ACaptureThresh[28]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[28]  ( .D(n7068), .CLK(n9214), .Q(
        ACaptureThresh_loc_reg_288[28]) );
  DFFPOSX1 \ACaptureThresh_reg[29]  ( .D(n4637), .CLK(n9214), .Q(
        ACaptureThresh[29]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[29]  ( .D(n7224), .CLK(n9214), .Q(
        ACaptureThresh_loc_reg_288[29]) );
  DFFPOSX1 \ACaptureThresh_reg[30]  ( .D(n4636), .CLK(n9213), .Q(
        ACaptureThresh[30]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[30]  ( .D(n7389), .CLK(n9213), .Q(
        ACaptureThresh_loc_reg_288[30]) );
  DFFPOSX1 \ACaptureThresh_reg[31]  ( .D(n4635), .CLK(n9213), .Q(
        ACaptureThresh[31]) );
  DFFPOSX1 \ACaptureThresh_loc_reg_288_reg[31]  ( .D(n7574), .CLK(n9213), .Q(
        ACaptureThresh_loc_reg_288[31]) );
  DFFPOSX1 \VCaptureThresh_reg[0]  ( .D(n4602), .CLK(n9213), .Q(
        VCaptureThresh[0]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[0]  ( .D(n7768), .CLK(n9213), .Q(
        VCaptureThresh_loc_reg_298[0]) );
  DFFPOSX1 \VCaptureThresh_reg[1]  ( .D(n4601), .CLK(n9213), .Q(
        VCaptureThresh[1]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[1]  ( .D(n8227), .CLK(n9213), .Q(
        VCaptureThresh_loc_reg_298[1]) );
  DFFPOSX1 \VCaptureThresh_reg[2]  ( .D(n4600), .CLK(n9213), .Q(
        VCaptureThresh[2]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[2]  ( .D(n6246), .CLK(n9213), .Q(
        VCaptureThresh_loc_reg_298[2]) );
  DFFPOSX1 \VCaptureThresh_reg[3]  ( .D(n4599), .CLK(n9213), .Q(
        VCaptureThresh[3]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[3]  ( .D(n6341), .CLK(n9213), .Q(
        VCaptureThresh_loc_reg_298[3]) );
  DFFPOSX1 \VCaptureThresh_reg[4]  ( .D(n4598), .CLK(n9213), .Q(
        VCaptureThresh[4]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[4]  ( .D(n6450), .CLK(n9212), .Q(
        VCaptureThresh_loc_reg_298[4]) );
  DFFPOSX1 \VCaptureThresh_reg[5]  ( .D(n4597), .CLK(n9212), .Q(
        VCaptureThresh[5]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[5]  ( .D(n6563), .CLK(n9212), .Q(
        VCaptureThresh_loc_reg_298[5]) );
  DFFPOSX1 \VCaptureThresh_reg[6]  ( .D(n4596), .CLK(n9212), .Q(
        VCaptureThresh[6]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[6]  ( .D(n7989), .CLK(n9212), .Q(
        VCaptureThresh_loc_reg_298[6]) );
  DFFPOSX1 \VCaptureThresh_reg[7]  ( .D(n4595), .CLK(n9212), .Q(
        VCaptureThresh[7]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[7]  ( .D(n6672), .CLK(n9212), .Q(
        VCaptureThresh_loc_reg_298[7]) );
  DFFPOSX1 \VCaptureThresh_reg[8]  ( .D(n4594), .CLK(n9212), .Q(
        VCaptureThresh[8]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[8]  ( .D(n6793), .CLK(n9212), .Q(
        VCaptureThresh_loc_reg_298[8]) );
  DFFPOSX1 \VCaptureThresh_reg[9]  ( .D(n4593), .CLK(n9212), .Q(
        VCaptureThresh[9]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[9]  ( .D(n6928), .CLK(n9212), .Q(
        VCaptureThresh_loc_reg_298[9]) );
  DFFPOSX1 \VCaptureThresh_reg[10]  ( .D(n4592), .CLK(n9212), .Q(
        VCaptureThresh[10]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[10]  ( .D(n7071), .CLK(n9212), .Q(
        VCaptureThresh_loc_reg_298[10]) );
  DFFPOSX1 \VCaptureThresh_reg[11]  ( .D(n4591), .CLK(n9211), .Q(
        VCaptureThresh[11]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[11]  ( .D(n7227), .CLK(n9211), .Q(
        VCaptureThresh_loc_reg_298[11]) );
  DFFPOSX1 \VCaptureThresh_reg[12]  ( .D(n4590), .CLK(n9211), .Q(
        VCaptureThresh[12]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[12]  ( .D(n7392), .CLK(n9211), .Q(
        VCaptureThresh_loc_reg_298[12]) );
  DFFPOSX1 \VCaptureThresh_reg[13]  ( .D(n4589), .CLK(n9211), .Q(
        VCaptureThresh[13]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[13]  ( .D(n7771), .CLK(n9211), .Q(
        VCaptureThresh_loc_reg_298[13]) );
  DFFPOSX1 \VCaptureThresh_reg[14]  ( .D(n4588), .CLK(n9211), .Q(
        VCaptureThresh[14]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[14]  ( .D(n8230), .CLK(n9211), .Q(
        VCaptureThresh_loc_reg_298[14]) );
  DFFPOSX1 \VCaptureThresh_reg[15]  ( .D(n4587), .CLK(n9211), .Q(
        VCaptureThresh[15]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[15]  ( .D(n7577), .CLK(n9211), .Q(
        VCaptureThresh_loc_reg_298[15]) );
  DFFPOSX1 \VCaptureThresh_reg[16]  ( .D(n4586), .CLK(n9211), .Q(
        VCaptureThresh[16]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[16]  ( .D(n6161), .CLK(n9211), .Q(
        VCaptureThresh_loc_reg_298[16]) );
  DFFPOSX1 \VCaptureThresh_reg[17]  ( .D(n4585), .CLK(n9211), .Q(
        VCaptureThresh[17]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[17]  ( .D(n6249), .CLK(n9210), .Q(
        VCaptureThresh_loc_reg_298[17]) );
  DFFPOSX1 \VCaptureThresh_reg[18]  ( .D(n4584), .CLK(n9210), .Q(
        VCaptureThresh[18]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[18]  ( .D(n6344), .CLK(n9210), .Q(
        VCaptureThresh_loc_reg_298[18]) );
  DFFPOSX1 \VCaptureThresh_reg[19]  ( .D(n4583), .CLK(n9210), .Q(
        VCaptureThresh[19]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[19]  ( .D(n7992), .CLK(n9210), .Q(
        VCaptureThresh_loc_reg_298[19]) );
  DFFPOSX1 \VCaptureThresh_reg[20]  ( .D(n4582), .CLK(n9210), .Q(
        VCaptureThresh[20]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[20]  ( .D(n6453), .CLK(n9210), .Q(
        VCaptureThresh_loc_reg_298[20]) );
  DFFPOSX1 \VCaptureThresh_reg[21]  ( .D(n4581), .CLK(n9210), .Q(
        VCaptureThresh[21]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[21]  ( .D(n6566), .CLK(n9210), .Q(
        VCaptureThresh_loc_reg_298[21]) );
  DFFPOSX1 \VCaptureThresh_reg[22]  ( .D(n4580), .CLK(n9210), .Q(
        VCaptureThresh[22]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[22]  ( .D(n6675), .CLK(n9210), .Q(
        VCaptureThresh_loc_reg_298[22]) );
  DFFPOSX1 \VCaptureThresh_reg[23]  ( .D(n4579), .CLK(n9210), .Q(
        VCaptureThresh[23]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[23]  ( .D(n6796), .CLK(n9210), .Q(
        VCaptureThresh_loc_reg_298[23]) );
  DFFPOSX1 \VCaptureThresh_reg[24]  ( .D(n4578), .CLK(n9209), .Q(
        VCaptureThresh[24]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[24]  ( .D(n6931), .CLK(n9209), .Q(
        VCaptureThresh_loc_reg_298[24]) );
  DFFPOSX1 \VCaptureThresh_reg[25]  ( .D(n4577), .CLK(n9209), .Q(
        VCaptureThresh[25]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[25]  ( .D(n7074), .CLK(n9209), .Q(
        VCaptureThresh_loc_reg_298[25]) );
  DFFPOSX1 \VCaptureThresh_reg[26]  ( .D(n4576), .CLK(n9209), .Q(
        VCaptureThresh[26]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[26]  ( .D(n7230), .CLK(n9209), .Q(
        VCaptureThresh_loc_reg_298[26]) );
  DFFPOSX1 \VCaptureThresh_reg[27]  ( .D(n4575), .CLK(n9209), .Q(
        VCaptureThresh[27]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[27]  ( .D(n7395), .CLK(n9209), .Q(
        VCaptureThresh_loc_reg_298[27]) );
  DFFPOSX1 \VCaptureThresh_reg[28]  ( .D(n4574), .CLK(n9209), .Q(
        VCaptureThresh[28]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[28]  ( .D(n7580), .CLK(n9209), .Q(
        VCaptureThresh_loc_reg_298[28]) );
  DFFPOSX1 \VCaptureThresh_reg[29]  ( .D(n4573), .CLK(n9209), .Q(
        VCaptureThresh[29]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[29]  ( .D(n7774), .CLK(n9209), .Q(
        VCaptureThresh_loc_reg_298[29]) );
  DFFPOSX1 \VCaptureThresh_reg[30]  ( .D(n4572), .CLK(n9209), .Q(
        VCaptureThresh[30]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[30]  ( .D(n8233), .CLK(n9208), .Q(
        VCaptureThresh_loc_reg_298[30]) );
  DFFPOSX1 \VCaptureThresh_reg[31]  ( .D(n4571), .CLK(n9208), .Q(
        VCaptureThresh[31]) );
  DFFPOSX1 \VCaptureThresh_loc_reg_298_reg[31]  ( .D(n7995), .CLK(n9208), .Q(
        VCaptureThresh_loc_reg_298[31]) );
  DFFPOSX1 \a_thresh_reg[0]  ( .D(n9434), .CLK(n9208), .Q(a_thresh[0]) );
  DFFPOSX1 \a_thresh_reg[1]  ( .D(n9435), .CLK(n9208), .Q(a_thresh[1]) );
  DFFPOSX1 \a_thresh_reg[2]  ( .D(n9436), .CLK(n9208), .Q(a_thresh[2]) );
  DFFPOSX1 \a_thresh_reg[3]  ( .D(n9437), .CLK(n9208), .Q(a_thresh[3]) );
  DFFPOSX1 \a_thresh_reg[4]  ( .D(n9438), .CLK(n9208), .Q(a_thresh[4]) );
  DFFPOSX1 \a_thresh_reg[5]  ( .D(n9439), .CLK(n9208), .Q(a_thresh[5]) );
  DFFPOSX1 \a_thresh_reg[6]  ( .D(n9440), .CLK(n9208), .Q(a_thresh[6]) );
  DFFPOSX1 \a_thresh_reg[7]  ( .D(n9441), .CLK(n9208), .Q(a_thresh[7]) );
  DFFPOSX1 \a_thresh_reg[8]  ( .D(n9442), .CLK(n9208), .Q(a_thresh[8]) );
  DFFPOSX1 \a_thresh_reg[9]  ( .D(n9443), .CLK(n9208), .Q(a_thresh[9]) );
  DFFPOSX1 \a_thresh_reg[10]  ( .D(n9444), .CLK(n9207), .Q(a_thresh[10]) );
  DFFPOSX1 \a_thresh_reg[11]  ( .D(n9445), .CLK(n9207), .Q(a_thresh[11]) );
  DFFPOSX1 \a_thresh_reg[12]  ( .D(n9446), .CLK(n9207), .Q(a_thresh[12]) );
  DFFPOSX1 \a_thresh_reg[13]  ( .D(n9447), .CLK(n9207), .Q(a_thresh[13]) );
  DFFPOSX1 \a_thresh_reg[14]  ( .D(n9448), .CLK(n9207), .Q(a_thresh[14]) );
  DFFPOSX1 \a_thresh_reg[15]  ( .D(n9449), .CLK(n9207), .Q(a_thresh[15]) );
  DFFPOSX1 \a_thresh_reg[16]  ( .D(n9450), .CLK(n9207), .Q(a_thresh[16]) );
  DFFPOSX1 \a_thresh_reg[17]  ( .D(n9451), .CLK(n9207), .Q(a_thresh[17]) );
  DFFPOSX1 \a_thresh_reg[18]  ( .D(n9452), .CLK(n9207), .Q(a_thresh[18]) );
  DFFPOSX1 \a_thresh_reg[19]  ( .D(n9453), .CLK(n9207), .Q(a_thresh[19]) );
  DFFPOSX1 \a_thresh_reg[20]  ( .D(n9454), .CLK(n9207), .Q(a_thresh[20]) );
  DFFPOSX1 \a_thresh_reg[21]  ( .D(n9455), .CLK(n9207), .Q(a_thresh[21]) );
  DFFPOSX1 \a_thresh_reg[22]  ( .D(n9456), .CLK(n9207), .Q(a_thresh[22]) );
  DFFPOSX1 \a_thresh_reg[23]  ( .D(n9457), .CLK(n9206), .Q(a_thresh[23]) );
  DFFPOSX1 \a_thresh_reg[24]  ( .D(n9458), .CLK(n9206), .Q(a_thresh[24]) );
  DFFPOSX1 \a_thresh_reg[25]  ( .D(n9459), .CLK(n9206), .Q(a_thresh[25]) );
  DFFPOSX1 \a_thresh_reg[26]  ( .D(n9460), .CLK(n9206), .Q(a_thresh[26]) );
  DFFPOSX1 \a_thresh_reg[27]  ( .D(n9461), .CLK(n9206), .Q(a_thresh[27]) );
  DFFPOSX1 \a_thresh_reg[28]  ( .D(n9462), .CLK(n9206), .Q(a_thresh[28]) );
  DFFPOSX1 \a_thresh_reg[29]  ( .D(n9463), .CLK(n9206), .Q(a_thresh[29]) );
  DFFPOSX1 \a_thresh_reg[30]  ( .D(n9464), .CLK(n9206), .Q(a_thresh[30]) );
  DFFPOSX1 \a_thresh_reg[31]  ( .D(n9465), .CLK(n9206), .Q(a_thresh[31]) );
  DFFPOSX1 \aflip_reg[0]  ( .D(n4538), .CLK(n9206), .Q(aflip[0]) );
  DFFPOSX1 \aflip_reg[1]  ( .D(n4537), .CLK(n9206), .Q(aflip[1]) );
  DFFPOSX1 \aflip_reg[2]  ( .D(n4536), .CLK(n9206), .Q(aflip[2]) );
  DFFPOSX1 \data_read_reg_1495_reg[15]  ( .D(n9401), .CLK(n9206), .Q(
        data_read_reg_1495[15]) );
  DFFPOSX1 \data_read_reg_1495_reg[14]  ( .D(n9400), .CLK(n9205), .Q(
        data_read_reg_1495[14]) );
  DFFPOSX1 \data_read_reg_1495_reg[13]  ( .D(n9399), .CLK(n9205), .Q(
        data_read_reg_1495[13]) );
  DFFPOSX1 \data_read_reg_1495_reg[12]  ( .D(n9398), .CLK(n9205), .Q(
        data_read_reg_1495[12]) );
  DFFPOSX1 \data_read_reg_1495_reg[11]  ( .D(n9397), .CLK(n9205), .Q(
        data_read_reg_1495[11]) );
  DFFPOSX1 \data_read_reg_1495_reg[10]  ( .D(n9396), .CLK(n9205), .Q(
        data_read_reg_1495[10]) );
  DFFPOSX1 \data_read_reg_1495_reg[9]  ( .D(n9395), .CLK(n9205), .Q(
        data_read_reg_1495[9]) );
  DFFPOSX1 \data_read_reg_1495_reg[8]  ( .D(n9394), .CLK(n9205), .Q(
        data_read_reg_1495[8]) );
  DFFPOSX1 \data_read_reg_1495_reg[7]  ( .D(n9393), .CLK(n9205), .Q(
        data_read_reg_1495[7]) );
  DFFPOSX1 \data_read_reg_1495_reg[6]  ( .D(n9392), .CLK(n9205), .Q(
        data_read_reg_1495[6]) );
  DFFPOSX1 \data_read_reg_1495_reg[5]  ( .D(n9391), .CLK(n9205), .Q(
        data_read_reg_1495[5]) );
  DFFPOSX1 \data_read_reg_1495_reg[4]  ( .D(n9390), .CLK(n9205), .Q(
        data_read_reg_1495[4]) );
  DFFPOSX1 \data_read_reg_1495_reg[3]  ( .D(n9389), .CLK(n9205), .Q(
        data_read_reg_1495[3]) );
  DFFPOSX1 \data_read_reg_1495_reg[2]  ( .D(n9388), .CLK(n9205), .Q(
        data_read_reg_1495[2]) );
  DFFPOSX1 \data_read_reg_1495_reg[1]  ( .D(n9387), .CLK(n9204), .Q(
        data_read_reg_1495[1]) );
  DFFPOSX1 \data_read_reg_1495_reg[0]  ( .D(n9386), .CLK(n9204), .Q(
        data_read_reg_1495[0]) );
  DFFPOSX1 \ap_CS_fsm_reg[1]  ( .D(N99), .CLK(n9204), .Q(ap_CS_fsm[1]) );
  DFFPOSX1 \recentdatapoints_len_reg[0]  ( .D(n4053), .CLK(n9204), .Q(
        recentdatapoints_len[0]) );
  DFFPOSX1 \recentdatapoints_len_reg[10]  ( .D(n4052), .CLK(n9204), .Q(
        recentdatapoints_len[10]) );
  DFFPOSX1 \recentdatapoints_len_reg[1]  ( .D(n4051), .CLK(n9204), .Q(
        recentdatapoints_len[1]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[1]  ( .D(n4050), .CLK(n9204), .Q(
        tmp_38_i_reg_1550[1]) );
  DFFPOSX1 \recentdatapoints_len_reg[2]  ( .D(n4049), .CLK(n9204), .Q(
        recentdatapoints_len[2]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[2]  ( .D(n4048), .CLK(n9204), .Q(
        tmp_38_i_reg_1550[2]) );
  DFFPOSX1 \recentdatapoints_len_reg[3]  ( .D(n4047), .CLK(n9204), .Q(
        recentdatapoints_len[3]) );
  DFFPOSX1 \recentdatapoints_len_reg[4]  ( .D(n4046), .CLK(n9204), .Q(
        recentdatapoints_len[4]) );
  DFFPOSX1 \recentdatapoints_len_reg[5]  ( .D(n4045), .CLK(n9204), .Q(
        recentdatapoints_len[5]) );
  DFFPOSX1 \recentdatapoints_len_reg[6]  ( .D(n4044), .CLK(n9204), .Q(
        recentdatapoints_len[6]) );
  DFFPOSX1 \recentdatapoints_len_reg[7]  ( .D(n4043), .CLK(n9203), .Q(
        recentdatapoints_len[7]) );
  DFFPOSX1 \recentdatapoints_len_reg[8]  ( .D(n4042), .CLK(n9203), .Q(
        recentdatapoints_len[8]) );
  DFFPOSX1 \recentdatapoints_len_reg[9]  ( .D(n4041), .CLK(n9203), .Q(
        recentdatapoints_len[9]) );
  DFFPOSX1 \recentdatapoints_len_reg[11]  ( .D(n4040), .CLK(n9203), .Q(
        recentdatapoints_len[11]) );
  DFFPOSX1 \recentdatapoints_len_reg[12]  ( .D(n4039), .CLK(n9203), .Q(
        recentdatapoints_len[12]) );
  DFFPOSX1 \recentdatapoints_len_reg[13]  ( .D(n4038), .CLK(n9203), .Q(
        recentdatapoints_len[13]) );
  DFFPOSX1 \recentdatapoints_len_reg[14]  ( .D(n4037), .CLK(n9203), .Q(
        recentdatapoints_len[14]) );
  DFFPOSX1 \recentdatapoints_len_reg[15]  ( .D(n4036), .CLK(n9203), .Q(
        recentdatapoints_len[15]) );
  DFFPOSX1 \recentdatapoints_len_reg[16]  ( .D(n4035), .CLK(n9203), .Q(
        recentdatapoints_len[16]) );
  DFFPOSX1 \recentdatapoints_len_reg[17]  ( .D(n4034), .CLK(n9203), .Q(
        recentdatapoints_len[17]) );
  DFFPOSX1 \recentdatapoints_len_reg[18]  ( .D(n4033), .CLK(n9203), .Q(
        recentdatapoints_len[18]) );
  DFFPOSX1 \recentdatapoints_len_reg[19]  ( .D(n4032), .CLK(n9203), .Q(
        recentdatapoints_len[19]) );
  DFFPOSX1 \recentdatapoints_len_reg[20]  ( .D(n4031), .CLK(n9203), .Q(
        recentdatapoints_len[20]) );
  DFFPOSX1 \recentdatapoints_len_reg[21]  ( .D(n4030), .CLK(n9202), .Q(
        recentdatapoints_len[21]) );
  DFFPOSX1 \recentdatapoints_len_reg[22]  ( .D(n4029), .CLK(n9202), .Q(
        recentdatapoints_len[22]) );
  DFFPOSX1 \recentdatapoints_len_reg[23]  ( .D(n4028), .CLK(n9202), .Q(
        recentdatapoints_len[23]) );
  DFFPOSX1 \recentdatapoints_len_reg[24]  ( .D(n4027), .CLK(n9202), .Q(
        recentdatapoints_len[24]) );
  DFFPOSX1 \recentdatapoints_len_reg[25]  ( .D(n4026), .CLK(n9202), .Q(
        recentdatapoints_len[25]) );
  DFFPOSX1 \recentdatapoints_len_reg[26]  ( .D(n4025), .CLK(n9202), .Q(
        recentdatapoints_len[26]) );
  DFFPOSX1 \recentdatapoints_len_reg[27]  ( .D(n4024), .CLK(n9202), .Q(
        recentdatapoints_len[27]) );
  DFFPOSX1 \recentdatapoints_len_reg[28]  ( .D(n4023), .CLK(n9202), .Q(
        recentdatapoints_len[28]) );
  DFFPOSX1 \recentdatapoints_len_reg[29]  ( .D(n4022), .CLK(n9202), .Q(
        recentdatapoints_len[29]) );
  DFFPOSX1 \recentdatapoints_len_reg[30]  ( .D(n4021), .CLK(n9202), .Q(
        recentdatapoints_len[30]) );
  DFFPOSX1 \recentdatapoints_len_reg[31]  ( .D(n4020), .CLK(n9202), .Q(
        recentdatapoints_len[31]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[0]  ( .D(n4019), .CLK(n9202), .Q(
        tmp_38_i_reg_1550[0]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[0]  ( .D(n4018), .CLK(n9202), .Q(
        recentdatapoints_head_i[0]) );
  DFFPOSX1 \recentdatapoints_data_addr_reg_1533_reg[0]  ( .D(n4017), .CLK(
        n9201), .Q(recentdatapoints_data_addr_reg_1533[0]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[1]  ( .D(n4016), .CLK(n9201), .Q(
        recentdatapoints_head_i[1]) );
  DFFPOSX1 \recentdatapoints_data_addr_reg_1533_reg[1]  ( .D(n4015), .CLK(
        n9201), .Q(recentdatapoints_data_addr_reg_1533[1]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[3]  ( .D(n4014), .CLK(n9201), .Q(
        recentdatapoints_head_i[3]) );
  DFFPOSX1 \recentdatapoints_data_addr_reg_1533_reg[3]  ( .D(n4013), .CLK(
        n9201), .Q(recentdatapoints_data_addr_reg_1533[3]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[5]  ( .D(n4012), .CLK(n9201), .Q(
        recentdatapoints_head_i[5]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[6]  ( .D(n4011), .CLK(n9201), .Q(
        recentdatapoints_head_i[6]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[7]  ( .D(n4010), .CLK(n9201), .Q(
        recentdatapoints_head_i[7]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[8]  ( .D(n4009), .CLK(n9201), .Q(
        recentdatapoints_head_i[8]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[9]  ( .D(n4008), .CLK(n9201), .Q(
        recentdatapoints_head_i[9]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[10]  ( .D(n4007), .CLK(n9201), .Q(
        recentdatapoints_head_i[10]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[11]  ( .D(n4006), .CLK(n9201), .Q(
        recentdatapoints_head_i[11]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[12]  ( .D(n4005), .CLK(n9201), .Q(
        recentdatapoints_head_i[12]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[13]  ( .D(n4004), .CLK(n9200), .Q(
        recentdatapoints_head_i[13]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[14]  ( .D(n4003), .CLK(n9200), .Q(
        recentdatapoints_head_i[14]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[15]  ( .D(n4002), .CLK(n9200), .Q(
        recentdatapoints_head_i[15]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[16]  ( .D(n4001), .CLK(n9200), .Q(
        recentdatapoints_head_i[16]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[17]  ( .D(n4000), .CLK(n9200), .Q(
        recentdatapoints_head_i[17]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[18]  ( .D(n3999), .CLK(n9200), .Q(
        recentdatapoints_head_i[18]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[19]  ( .D(n3998), .CLK(n9200), .Q(
        recentdatapoints_head_i[19]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[20]  ( .D(n3997), .CLK(n9200), .Q(
        recentdatapoints_head_i[20]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[21]  ( .D(n3996), .CLK(n9200), .Q(
        recentdatapoints_head_i[21]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[22]  ( .D(n3995), .CLK(n9200), .Q(
        recentdatapoints_head_i[22]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[23]  ( .D(n3994), .CLK(n9200), .Q(
        recentdatapoints_head_i[23]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[24]  ( .D(n3993), .CLK(n9200), .Q(
        recentdatapoints_head_i[24]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[25]  ( .D(n3992), .CLK(n9200), .Q(
        recentdatapoints_head_i[25]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[26]  ( .D(n3991), .CLK(n9199), .Q(
        recentdatapoints_head_i[26]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[27]  ( .D(n3990), .CLK(n9199), .Q(
        recentdatapoints_head_i[27]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[28]  ( .D(n3989), .CLK(n9199), .Q(
        recentdatapoints_head_i[28]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[29]  ( .D(n3988), .CLK(n9199), .Q(
        recentdatapoints_head_i[29]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[30]  ( .D(n3987), .CLK(n9199), .Q(
        recentdatapoints_head_i[30]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[31]  ( .D(n3986), .CLK(n9199), .Q(
        recentdatapoints_head_i[31]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[4]  ( .D(n3985), .CLK(n9199), .Q(
        recentdatapoints_head_i[4]) );
  DFFPOSX1 \recentdatapoints_data_addr_reg_1533_reg[4]  ( .D(n3984), .CLK(
        n9199), .Q(recentdatapoints_data_addr_reg_1533[4]) );
  DFFPOSX1 \recentdatapoints_head_i_reg[2]  ( .D(n3983), .CLK(n9199), .Q(
        recentdatapoints_head_i[2]) );
  DFFPOSX1 \recentdatapoints_data_addr_reg_1533_reg[2]  ( .D(n3982), .CLK(
        n9199), .Q(recentdatapoints_data_addr_reg_1533[2]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[31]  ( .D(n3981), .CLK(n9199), .Q(
        p_tmp_i_reg_1556[31]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[30]  ( .D(n3980), .CLK(n9199), .Q(
        p_tmp_i_reg_1556[30]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[29]  ( .D(n3979), .CLK(n9199), .Q(
        p_tmp_i_reg_1556[29]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[28]  ( .D(n3978), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[28]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[27]  ( .D(n3977), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[27]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[26]  ( .D(n3976), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[26]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[25]  ( .D(n3975), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[25]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[24]  ( .D(n3974), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[24]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[23]  ( .D(n3973), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[23]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[22]  ( .D(n3972), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[22]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[21]  ( .D(n3971), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[21]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[20]  ( .D(n3970), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[20]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[19]  ( .D(n3969), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[19]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[18]  ( .D(n3968), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[18]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[17]  ( .D(n3967), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[17]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[16]  ( .D(n3966), .CLK(n9198), .Q(
        p_tmp_i_reg_1556[16]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[15]  ( .D(n3965), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[15]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[14]  ( .D(n3964), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[14]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[13]  ( .D(n3963), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[13]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[12]  ( .D(n3962), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[12]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[11]  ( .D(n3961), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[11]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[10]  ( .D(n3960), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[10]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[9]  ( .D(n3959), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[9]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[8]  ( .D(n3958), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[8]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[7]  ( .D(n3957), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[7]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[6]  ( .D(n3956), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[6]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[5]  ( .D(n3955), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[5]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[4]  ( .D(n3954), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[4]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[3]  ( .D(n3953), .CLK(n9197), .Q(
        p_tmp_i_reg_1556[3]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[2]  ( .D(n3952), .CLK(n9196), .Q(
        p_tmp_i_reg_1556[2]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[1]  ( .D(n3951), .CLK(n9196), .Q(
        p_tmp_i_reg_1556[1]) );
  DFFPOSX1 \p_tmp_i_reg_1556_reg[0]  ( .D(n3950), .CLK(n9196), .Q(
        p_tmp_i_reg_1556[0]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[31]  ( .D(n3949), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[31]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[30]  ( .D(n3948), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[30]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[29]  ( .D(n3947), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[29]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[28]  ( .D(n3946), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[28]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[27]  ( .D(n3945), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[27]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[26]  ( .D(n3944), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[26]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[25]  ( .D(n3943), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[25]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[24]  ( .D(n3942), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[24]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[23]  ( .D(n3941), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[23]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[22]  ( .D(n3940), .CLK(n9196), .Q(
        tmp_38_i_reg_1550[22]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[21]  ( .D(n3939), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[21]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[20]  ( .D(n3938), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[20]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[19]  ( .D(n3937), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[19]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[18]  ( .D(n3936), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[18]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[17]  ( .D(n3935), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[17]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[16]  ( .D(n3934), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[16]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[15]  ( .D(n3933), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[15]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[14]  ( .D(n3932), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[14]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[13]  ( .D(n3931), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[13]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[12]  ( .D(n3930), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[12]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[11]  ( .D(n3929), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[11]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[10]  ( .D(n3928), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[10]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[9]  ( .D(n3927), .CLK(n9195), .Q(
        tmp_38_i_reg_1550[9]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[8]  ( .D(n3926), .CLK(n9194), .Q(
        tmp_38_i_reg_1550[8]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[7]  ( .D(n3925), .CLK(n9194), .Q(
        tmp_38_i_reg_1550[7]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[6]  ( .D(n3924), .CLK(n9194), .Q(
        tmp_38_i_reg_1550[6]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[5]  ( .D(n3923), .CLK(n9194), .Q(
        tmp_38_i_reg_1550[5]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[4]  ( .D(n3922), .CLK(n9194), .Q(
        tmp_38_i_reg_1550[4]) );
  DFFPOSX1 \tmp_38_i_reg_1550_reg[3]  ( .D(n3921), .CLK(n9194), .Q(
        tmp_38_i_reg_1550[3]) );
  DFFPOSX1 \ap_CS_fsm_reg[2]  ( .D(N100), .CLK(n9194), .Q(ap_CS_fsm[2]) );
  DFFPOSX1 \ap_CS_fsm_reg[3]  ( .D(N101), .CLK(n9194), .Q(ap_CS_fsm[3]) );
  DFFPOSX1 \ap_CS_fsm_reg[4]  ( .D(N102), .CLK(n9194), .Q(ap_CS_fsm[4]) );
  DFFPOSX1 \recentVBools_head_i_reg[3]  ( .D(n3920), .CLK(n9194), .Q(
        recentVBools_head_i[3]) );
  DFFPOSX1 \recentVBools_data_addr_reg_1573_reg[3]  ( .D(n3919), .CLK(n9194), 
        .Q(recentVBools_data_addr_reg_1573[3]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[0]  ( .D(n3918), .CLK(
        n9194), .Q(CircularBuffer_head_i_read_ass_reg_1624[0]) );
  DFFPOSX1 \recentVBools_head_i_reg[0]  ( .D(n3917), .CLK(n9194), .Q(
        recentVBools_head_i[0]) );
  DFFPOSX1 \recentVBools_data_addr_reg_1573_reg[0]  ( .D(n3916), .CLK(n9193), 
        .Q(recentVBools_data_addr_reg_1573[0]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[5]  ( .D(n3915), .CLK(
        n9193), .Q(CircularBuffer_head_i_read_ass_reg_1624[5]) );
  DFFPOSX1 \recentVBools_head_i_reg[5]  ( .D(n3914), .CLK(n9193), .Q(
        recentVBools_head_i[5]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[6]  ( .D(n3913), .CLK(
        n9193), .Q(CircularBuffer_head_i_read_ass_reg_1624[6]) );
  DFFPOSX1 \recentVBools_head_i_reg[6]  ( .D(n3912), .CLK(n9193), .Q(
        recentVBools_head_i[6]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[7]  ( .D(n3911), .CLK(
        n9193), .Q(CircularBuffer_head_i_read_ass_reg_1624[7]) );
  DFFPOSX1 \recentVBools_head_i_reg[7]  ( .D(n3910), .CLK(n9193), .Q(
        recentVBools_head_i[7]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[8]  ( .D(n3909), .CLK(
        n9193), .Q(CircularBuffer_head_i_read_ass_reg_1624[8]) );
  DFFPOSX1 \recentVBools_head_i_reg[8]  ( .D(n3908), .CLK(n9193), .Q(
        recentVBools_head_i[8]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[9]  ( .D(n3907), .CLK(
        n9193), .Q(CircularBuffer_head_i_read_ass_reg_1624[9]) );
  DFFPOSX1 \recentVBools_head_i_reg[9]  ( .D(n3906), .CLK(n9193), .Q(
        recentVBools_head_i[9]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[10]  ( .D(n3905), 
        .CLK(n9193), .Q(CircularBuffer_head_i_read_ass_reg_1624[10]) );
  DFFPOSX1 \recentVBools_head_i_reg[10]  ( .D(n3904), .CLK(n9193), .Q(
        recentVBools_head_i[10]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[11]  ( .D(n3903), 
        .CLK(n9192), .Q(CircularBuffer_head_i_read_ass_reg_1624[11]) );
  DFFPOSX1 \recentVBools_head_i_reg[11]  ( .D(n3902), .CLK(n9192), .Q(
        recentVBools_head_i[11]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[12]  ( .D(n3901), 
        .CLK(n9192), .Q(CircularBuffer_head_i_read_ass_reg_1624[12]) );
  DFFPOSX1 \recentVBools_head_i_reg[12]  ( .D(n3900), .CLK(n9192), .Q(
        recentVBools_head_i[12]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[13]  ( .D(n3899), 
        .CLK(n9192), .Q(CircularBuffer_head_i_read_ass_reg_1624[13]) );
  DFFPOSX1 \recentVBools_head_i_reg[13]  ( .D(n3898), .CLK(n9192), .Q(
        recentVBools_head_i[13]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[14]  ( .D(n3897), 
        .CLK(n9192), .Q(CircularBuffer_head_i_read_ass_reg_1624[14]) );
  DFFPOSX1 \recentVBools_head_i_reg[14]  ( .D(n3896), .CLK(n9192), .Q(
        recentVBools_head_i[14]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[15]  ( .D(n3895), 
        .CLK(n9192), .Q(CircularBuffer_head_i_read_ass_reg_1624[15]) );
  DFFPOSX1 \recentVBools_head_i_reg[15]  ( .D(n3894), .CLK(n9192), .Q(
        recentVBools_head_i[15]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[16]  ( .D(n3893), 
        .CLK(n9192), .Q(CircularBuffer_head_i_read_ass_reg_1624[16]) );
  DFFPOSX1 \recentVBools_head_i_reg[16]  ( .D(n3892), .CLK(n9192), .Q(
        recentVBools_head_i[16]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[17]  ( .D(n3891), 
        .CLK(n9192), .Q(CircularBuffer_head_i_read_ass_reg_1624[17]) );
  DFFPOSX1 \recentVBools_head_i_reg[17]  ( .D(n3890), .CLK(n9191), .Q(
        recentVBools_head_i[17]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[18]  ( .D(n3889), 
        .CLK(n9191), .Q(CircularBuffer_head_i_read_ass_reg_1624[18]) );
  DFFPOSX1 \recentVBools_head_i_reg[18]  ( .D(n3888), .CLK(n9191), .Q(
        recentVBools_head_i[18]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[19]  ( .D(n3887), 
        .CLK(n9191), .Q(CircularBuffer_head_i_read_ass_reg_1624[19]) );
  DFFPOSX1 \recentVBools_head_i_reg[19]  ( .D(n3886), .CLK(n9191), .Q(
        recentVBools_head_i[19]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[20]  ( .D(n3885), 
        .CLK(n9191), .Q(CircularBuffer_head_i_read_ass_reg_1624[20]) );
  DFFPOSX1 \recentVBools_head_i_reg[20]  ( .D(n3884), .CLK(n9191), .Q(
        recentVBools_head_i[20]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[21]  ( .D(n3883), 
        .CLK(n9191), .Q(CircularBuffer_head_i_read_ass_reg_1624[21]) );
  DFFPOSX1 \recentVBools_head_i_reg[21]  ( .D(n3882), .CLK(n9191), .Q(
        recentVBools_head_i[21]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[22]  ( .D(n3881), 
        .CLK(n9191), .Q(CircularBuffer_head_i_read_ass_reg_1624[22]) );
  DFFPOSX1 \recentVBools_head_i_reg[22]  ( .D(n3880), .CLK(n9191), .Q(
        recentVBools_head_i[22]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[23]  ( .D(n3879), 
        .CLK(n9191), .Q(CircularBuffer_head_i_read_ass_reg_1624[23]) );
  DFFPOSX1 \recentVBools_head_i_reg[23]  ( .D(n3878), .CLK(n9191), .Q(
        recentVBools_head_i[23]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[24]  ( .D(n3877), 
        .CLK(n9190), .Q(CircularBuffer_head_i_read_ass_reg_1624[24]) );
  DFFPOSX1 \recentVBools_head_i_reg[24]  ( .D(n3876), .CLK(n9190), .Q(
        recentVBools_head_i[24]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[25]  ( .D(n3875), 
        .CLK(n9190), .Q(CircularBuffer_head_i_read_ass_reg_1624[25]) );
  DFFPOSX1 \recentVBools_head_i_reg[25]  ( .D(n3874), .CLK(n9190), .Q(
        recentVBools_head_i[25]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[26]  ( .D(n3873), 
        .CLK(n9190), .Q(CircularBuffer_head_i_read_ass_reg_1624[26]) );
  DFFPOSX1 \recentVBools_head_i_reg[26]  ( .D(n3872), .CLK(n9190), .Q(
        recentVBools_head_i[26]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[27]  ( .D(n3871), 
        .CLK(n9190), .Q(CircularBuffer_head_i_read_ass_reg_1624[27]) );
  DFFPOSX1 \recentVBools_head_i_reg[27]  ( .D(n3870), .CLK(n9190), .Q(
        recentVBools_head_i[27]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[28]  ( .D(n3869), 
        .CLK(n9190), .Q(CircularBuffer_head_i_read_ass_reg_1624[28]) );
  DFFPOSX1 \recentVBools_head_i_reg[28]  ( .D(n3868), .CLK(n9190), .Q(
        recentVBools_head_i[28]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[29]  ( .D(n3867), 
        .CLK(n9190), .Q(CircularBuffer_head_i_read_ass_reg_1624[29]) );
  DFFPOSX1 \recentVBools_head_i_reg[29]  ( .D(n3866), .CLK(n9190), .Q(
        recentVBools_head_i[29]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[30]  ( .D(n3865), 
        .CLK(n9190), .Q(CircularBuffer_head_i_read_ass_reg_1624[30]) );
  DFFPOSX1 \recentVBools_head_i_reg[30]  ( .D(n3864), .CLK(n9189), .Q(
        recentVBools_head_i[30]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[31]  ( .D(n3863), 
        .CLK(n9189), .Q(CircularBuffer_head_i_read_ass_reg_1624[31]) );
  DFFPOSX1 \recentVBools_head_i_reg[31]  ( .D(n3862), .CLK(n9189), .Q(
        recentVBools_head_i[31]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[4]  ( .D(n7563), .CLK(
        n9189), .Q(CircularBuffer_head_i_read_ass_reg_1624[4]) );
  DFFPOSX1 \recentVBools_head_i_reg[4]  ( .D(n3860), .CLK(n9189), .Q(
        recentVBools_head_i[4]) );
  DFFPOSX1 \recentVBools_data_addr_reg_1573_reg[4]  ( .D(n3859), .CLK(n9189), 
        .Q(recentVBools_data_addr_reg_1573[4]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[3]  ( .D(n7382), .CLK(
        n9189), .Q(CircularBuffer_head_i_read_ass_reg_1624[3]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[2]  ( .D(n7761), .CLK(
        n9189), .Q(CircularBuffer_head_i_read_ass_reg_1624[2]) );
  DFFPOSX1 \recentVBools_head_i_reg[2]  ( .D(n3856), .CLK(n9189), .Q(
        recentVBools_head_i[2]) );
  DFFPOSX1 \recentVBools_data_addr_reg_1573_reg[2]  ( .D(n3855), .CLK(n9189), 
        .Q(recentVBools_data_addr_reg_1573[2]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_reg_1624_reg[1]  ( .D(n7979), .CLK(
        n9189), .Q(CircularBuffer_head_i_read_ass_reg_1624[1]) );
  DFFPOSX1 \recentVBools_head_i_reg[1]  ( .D(n3853), .CLK(n9189), .Q(
        recentVBools_head_i[1]) );
  DFFPOSX1 \recentVBools_data_addr_reg_1573_reg[1]  ( .D(n3852), .CLK(n9189), 
        .Q(recentVBools_data_addr_reg_1573[1]) );
  DFFPOSX1 \ap_CS_fsm_reg[5]  ( .D(N103), .CLK(n9188), .Q(ap_CS_fsm[5]) );
  DFFPOSX1 \ap_CS_fsm_reg[6]  ( .D(N104), .CLK(n9188), .Q(ap_CS_fsm[6]) );
  DFFPOSX1 \ap_CS_fsm_reg[7]  ( .D(n4759), .CLK(n9188), .Q(ap_CS_fsm[7]) );
  DFFPOSX1 \tmp_i3_reg_1674_reg[0]  ( .D(n3851), .CLK(n9188), .Q(
        \tmp_i3_reg_1674[0] ) );
  DFFPOSX1 \recentVBools_len_reg[0]  ( .D(n4534), .CLK(n9188), .Q(
        recentVBools_len[0]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[0]  ( .D(n3850), 
        .CLK(n9188), .Q(CircularBuffer_len_write_assig_1_fu_924_p2[0]) );
  DFFPOSX1 \tmp_8_reg_1630_reg[0]  ( .D(n3849), .CLK(n9188), .Q(
        \tmp_8_reg_1630[0] ) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[30]  ( .D(n4472), .CLK(n9188), 
        .Q(recentVBools_len_new_reg_317[30]) );
  DFFPOSX1 \recentVBools_len_reg[30]  ( .D(n4504), .CLK(n9188), .Q(
        recentVBools_len[30]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[1]  ( .D(n3848), 
        .CLK(n9188), .Q(CircularBuffer_len_read_assign_1_reg_1616[1]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[2]  ( .D(n3847), 
        .CLK(n9188), .Q(CircularBuffer_len_read_assign_1_reg_1616[2]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[3]  ( .D(n3846), 
        .CLK(n9188), .Q(CircularBuffer_len_read_assign_1_reg_1616[3]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[4]  ( .D(n3845), 
        .CLK(n9188), .Q(CircularBuffer_len_read_assign_1_reg_1616[4]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[5]  ( .D(n3844), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[5]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[6]  ( .D(n3843), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[6]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[7]  ( .D(n3842), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[7]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[8]  ( .D(n3841), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[8]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[9]  ( .D(n3840), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[9]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[10]  ( .D(n3839), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[10]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[11]  ( .D(n3838), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[11]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[12]  ( .D(n3837), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[12]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[13]  ( .D(n3836), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[13]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[14]  ( .D(n3835), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[14]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[15]  ( .D(n3834), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[15]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[16]  ( .D(n3833), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[16]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[17]  ( .D(n3832), 
        .CLK(n9187), .Q(CircularBuffer_len_read_assign_1_reg_1616[17]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[18]  ( .D(n3831), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[18]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[19]  ( .D(n3830), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[19]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[20]  ( .D(n3829), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[20]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[21]  ( .D(n3828), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[21]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[22]  ( .D(n3827), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[22]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[23]  ( .D(n3826), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[23]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[24]  ( .D(n3825), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[24]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[25]  ( .D(n3824), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[25]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[26]  ( .D(n3823), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[26]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[27]  ( .D(n3822), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[27]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[28]  ( .D(n3821), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[28]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[29]  ( .D(n3820), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[29]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[30]  ( .D(n3819), 
        .CLK(n9186), .Q(CircularBuffer_len_read_assign_1_reg_1616[30]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_1_reg_1616_reg[31]  ( .D(n3818), 
        .CLK(n9185), .Q(CircularBuffer_len_read_assign_1_reg_1616[31]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[1]  ( .D(n4501), .CLK(n9185), .Q(
        recentVBools_len_new_reg_317[1]) );
  DFFPOSX1 \recentVBools_len_reg[1]  ( .D(n4533), .CLK(n9185), .Q(
        recentVBools_len[1]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[2]  ( .D(n4500), .CLK(n9185), .Q(
        recentVBools_len_new_reg_317[2]) );
  DFFPOSX1 \recentVBools_len_reg[2]  ( .D(n4532), .CLK(n9185), .Q(
        recentVBools_len[2]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[3]  ( .D(n4499), .CLK(n9185), .Q(
        recentVBools_len_new_reg_317[3]) );
  DFFPOSX1 \recentVBools_len_reg[3]  ( .D(n4531), .CLK(n9185), .Q(
        recentVBools_len[3]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[4]  ( .D(n4498), .CLK(n9185), .Q(
        recentVBools_len_new_reg_317[4]) );
  DFFPOSX1 \recentVBools_len_reg[4]  ( .D(n4530), .CLK(n9185), .Q(
        recentVBools_len[4]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[5]  ( .D(n4497), .CLK(n9185), .Q(
        recentVBools_len_new_reg_317[5]) );
  DFFPOSX1 \recentVBools_len_reg[5]  ( .D(n4529), .CLK(n9185), .Q(
        recentVBools_len[5]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[6]  ( .D(n4496), .CLK(n9185), .Q(
        recentVBools_len_new_reg_317[6]) );
  DFFPOSX1 \recentVBools_len_reg[6]  ( .D(n4528), .CLK(n9185), .Q(
        recentVBools_len[6]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[7]  ( .D(n4495), .CLK(n9184), .Q(
        recentVBools_len_new_reg_317[7]) );
  DFFPOSX1 \recentVBools_len_reg[7]  ( .D(n4527), .CLK(n9184), .Q(
        recentVBools_len[7]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[8]  ( .D(n4494), .CLK(n9184), .Q(
        recentVBools_len_new_reg_317[8]) );
  DFFPOSX1 \recentVBools_len_reg[8]  ( .D(n4526), .CLK(n9184), .Q(
        recentVBools_len[8]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[9]  ( .D(n4493), .CLK(n9184), .Q(
        recentVBools_len_new_reg_317[9]) );
  DFFPOSX1 \recentVBools_len_reg[9]  ( .D(n4525), .CLK(n9184), .Q(
        recentVBools_len[9]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[10]  ( .D(n4492), .CLK(n9184), 
        .Q(recentVBools_len_new_reg_317[10]) );
  DFFPOSX1 \recentVBools_len_reg[10]  ( .D(n4524), .CLK(n9184), .Q(
        recentVBools_len[10]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[11]  ( .D(n4491), .CLK(n9184), 
        .Q(recentVBools_len_new_reg_317[11]) );
  DFFPOSX1 \recentVBools_len_reg[11]  ( .D(n4523), .CLK(n9184), .Q(
        recentVBools_len[11]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[12]  ( .D(n4490), .CLK(n9184), 
        .Q(recentVBools_len_new_reg_317[12]) );
  DFFPOSX1 \recentVBools_len_reg[12]  ( .D(n4522), .CLK(n9184), .Q(
        recentVBools_len[12]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[13]  ( .D(n4489), .CLK(n9184), 
        .Q(recentVBools_len_new_reg_317[13]) );
  DFFPOSX1 \recentVBools_len_reg[13]  ( .D(n4521), .CLK(n9183), .Q(
        recentVBools_len[13]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[14]  ( .D(n4488), .CLK(n9183), 
        .Q(recentVBools_len_new_reg_317[14]) );
  DFFPOSX1 \recentVBools_len_reg[14]  ( .D(n4520), .CLK(n9183), .Q(
        recentVBools_len[14]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[15]  ( .D(n4487), .CLK(n9183), 
        .Q(recentVBools_len_new_reg_317[15]) );
  DFFPOSX1 \recentVBools_len_reg[15]  ( .D(n4519), .CLK(n9183), .Q(
        recentVBools_len[15]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[16]  ( .D(n4486), .CLK(n9183), 
        .Q(recentVBools_len_new_reg_317[16]) );
  DFFPOSX1 \recentVBools_len_reg[16]  ( .D(n4518), .CLK(n9183), .Q(
        recentVBools_len[16]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[17]  ( .D(n4485), .CLK(n9183), 
        .Q(recentVBools_len_new_reg_317[17]) );
  DFFPOSX1 \recentVBools_len_reg[17]  ( .D(n4517), .CLK(n9183), .Q(
        recentVBools_len[17]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[18]  ( .D(n4484), .CLK(n9183), 
        .Q(recentVBools_len_new_reg_317[18]) );
  DFFPOSX1 \recentVBools_len_reg[18]  ( .D(n4516), .CLK(n9183), .Q(
        recentVBools_len[18]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[19]  ( .D(n4483), .CLK(n9183), 
        .Q(recentVBools_len_new_reg_317[19]) );
  DFFPOSX1 \recentVBools_len_reg[19]  ( .D(n4515), .CLK(n9183), .Q(
        recentVBools_len[19]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[20]  ( .D(n4482), .CLK(n9182), 
        .Q(recentVBools_len_new_reg_317[20]) );
  DFFPOSX1 \recentVBools_len_reg[20]  ( .D(n4514), .CLK(n9182), .Q(
        recentVBools_len[20]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[21]  ( .D(n4481), .CLK(n9182), 
        .Q(recentVBools_len_new_reg_317[21]) );
  DFFPOSX1 \recentVBools_len_reg[21]  ( .D(n4513), .CLK(n9182), .Q(
        recentVBools_len[21]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[22]  ( .D(n4480), .CLK(n9182), 
        .Q(recentVBools_len_new_reg_317[22]) );
  DFFPOSX1 \recentVBools_len_reg[22]  ( .D(n4512), .CLK(n9182), .Q(
        recentVBools_len[22]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[23]  ( .D(n4479), .CLK(n9182), 
        .Q(recentVBools_len_new_reg_317[23]) );
  DFFPOSX1 \recentVBools_len_reg[23]  ( .D(n4511), .CLK(n9182), .Q(
        recentVBools_len[23]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[24]  ( .D(n4478), .CLK(n9182), 
        .Q(recentVBools_len_new_reg_317[24]) );
  DFFPOSX1 \recentVBools_len_reg[24]  ( .D(n4510), .CLK(n9182), .Q(
        recentVBools_len[24]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[25]  ( .D(n4477), .CLK(n9182), 
        .Q(recentVBools_len_new_reg_317[25]) );
  DFFPOSX1 \recentVBools_len_reg[25]  ( .D(n4509), .CLK(n9182), .Q(
        recentVBools_len[25]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[26]  ( .D(n4476), .CLK(n9182), 
        .Q(recentVBools_len_new_reg_317[26]) );
  DFFPOSX1 \recentVBools_len_reg[26]  ( .D(n4508), .CLK(n9181), .Q(
        recentVBools_len[26]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[27]  ( .D(n4475), .CLK(n9181), 
        .Q(recentVBools_len_new_reg_317[27]) );
  DFFPOSX1 \recentVBools_len_reg[27]  ( .D(n4507), .CLK(n9181), .Q(
        recentVBools_len[27]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[28]  ( .D(n4474), .CLK(n9181), 
        .Q(recentVBools_len_new_reg_317[28]) );
  DFFPOSX1 \recentVBools_len_reg[28]  ( .D(n4506), .CLK(n9181), .Q(
        recentVBools_len[28]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[29]  ( .D(n4473), .CLK(n9181), 
        .Q(recentVBools_len_new_reg_317[29]) );
  DFFPOSX1 \recentVBools_len_reg[29]  ( .D(n4505), .CLK(n9181), .Q(
        recentVBools_len[29]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[0]  ( .D(n3817), .CLK(
        n9181), .Q(CircularBuffer_len_write_assig_reg_1634[0]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[1]  ( .D(n3816), .CLK(
        n9181), .Q(CircularBuffer_len_write_assig_reg_1634[1]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[2]  ( .D(n3815), .CLK(
        n9181), .Q(CircularBuffer_len_write_assig_reg_1634[2]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[3]  ( .D(n3814), .CLK(
        n9181), .Q(CircularBuffer_len_write_assig_reg_1634[3]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[4]  ( .D(n3813), .CLK(
        n9181), .Q(CircularBuffer_len_write_assig_reg_1634[4]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[5]  ( .D(n3812), .CLK(
        n9181), .Q(CircularBuffer_len_write_assig_reg_1634[5]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[6]  ( .D(n3811), .CLK(
        n9180), .Q(CircularBuffer_len_write_assig_reg_1634[6]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[7]  ( .D(n3810), .CLK(
        n9180), .Q(CircularBuffer_len_write_assig_reg_1634[7]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[8]  ( .D(n3809), .CLK(
        n9180), .Q(CircularBuffer_len_write_assig_reg_1634[8]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[9]  ( .D(n3808), .CLK(
        n9180), .Q(CircularBuffer_len_write_assig_reg_1634[9]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[10]  ( .D(n3807), 
        .CLK(n9180), .Q(CircularBuffer_len_write_assig_reg_1634[10]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[11]  ( .D(n3806), 
        .CLK(n9180), .Q(CircularBuffer_len_write_assig_reg_1634[11]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[12]  ( .D(n3805), 
        .CLK(n9180), .Q(CircularBuffer_len_write_assig_reg_1634[12]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[13]  ( .D(n3804), 
        .CLK(n9180), .Q(CircularBuffer_len_write_assig_reg_1634[13]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[14]  ( .D(n3803), 
        .CLK(n9180), .Q(CircularBuffer_len_write_assig_reg_1634[14]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[15]  ( .D(n3802), 
        .CLK(n9180), .Q(CircularBuffer_len_write_assig_reg_1634[15]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[16]  ( .D(n3801), 
        .CLK(n9180), .Q(CircularBuffer_len_write_assig_reg_1634[16]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[17]  ( .D(n3800), 
        .CLK(n9180), .Q(CircularBuffer_len_write_assig_reg_1634[17]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[18]  ( .D(n3799), 
        .CLK(n9180), .Q(CircularBuffer_len_write_assig_reg_1634[18]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[19]  ( .D(n3798), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[19]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[20]  ( .D(n3797), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[20]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[21]  ( .D(n3796), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[21]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[22]  ( .D(n3795), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[22]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[23]  ( .D(n3794), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[23]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[24]  ( .D(n3793), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[24]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[25]  ( .D(n3792), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[25]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[26]  ( .D(n3791), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[26]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[27]  ( .D(n3790), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[27]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[28]  ( .D(n3789), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[28]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[29]  ( .D(n3788), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[29]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[30]  ( .D(n3787), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[30]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_reg_1634_reg[31]  ( .D(n3786), 
        .CLK(n9179), .Q(CircularBuffer_len_write_assig_reg_1634[31]) );
  DFFPOSX1 \not_tmp_i_i4_reg_1650_reg[0]  ( .D(n4716), .CLK(n9178), .Q(
        \not_tmp_i_i4_reg_1650[0] ) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[31]  ( .D(n4535), .CLK(n9178), 
        .Q(recentVBools_len_new_reg_317[31]) );
  DFFPOSX1 \recentVBools_len_reg[31]  ( .D(n4503), .CLK(n9178), .Q(
        recentVBools_len[31]) );
  DFFPOSX1 \recentVBools_len_new_reg_317_reg[0]  ( .D(n4502), .CLK(n9178), .Q(
        recentVBools_len_new_reg_317[0]) );
  DFFPOSX1 \tmp_s_reg_1578_reg[0]  ( .D(n9496), .CLK(n9178), .Q(
        \tmp_s_reg_1578[0] ) );
  DFFPOSX1 \toReturn_6_reg_1660_reg[0]  ( .D(n8221), .CLK(n9178), .Q(
        \toReturn_6_reg_1660[0] ) );
  DFFPOSX1 \recentVBools_data_load_reg_1584_reg[0]  ( .D(n3782), .CLK(n9178), 
        .Q(\recentVBools_data_load_reg_1584[0] ) );
  DFFPOSX1 \toReturn_5_reg_1655_reg[0]  ( .D(n3781), .CLK(n9178), .Q(
        \toReturn_5_reg_1655[0] ) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[0]  ( .D(n3780), .CLK(
        n9178), .Q(CircularBuffer_sum_read_assign_reg_1610[0]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[1]  ( .D(n3779), .CLK(
        n9178), .Q(CircularBuffer_sum_read_assign_reg_1610[1]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[2]  ( .D(n3778), .CLK(
        n9178), .Q(CircularBuffer_sum_read_assign_reg_1610[2]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[3]  ( .D(n3777), .CLK(
        n9178), .Q(CircularBuffer_sum_read_assign_reg_1610[3]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[4]  ( .D(n3776), .CLK(
        n9178), .Q(CircularBuffer_sum_read_assign_reg_1610[4]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[5]  ( .D(n3775), .CLK(
        n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[5]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[6]  ( .D(n3774), .CLK(
        n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[6]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[7]  ( .D(n3773), .CLK(
        n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[7]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[8]  ( .D(n3772), .CLK(
        n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[8]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[9]  ( .D(n3771), .CLK(
        n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[9]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[10]  ( .D(n3770), 
        .CLK(n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[10]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[11]  ( .D(n3769), 
        .CLK(n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[11]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[12]  ( .D(n3768), 
        .CLK(n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[12]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[13]  ( .D(n3767), 
        .CLK(n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[13]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[14]  ( .D(n3766), 
        .CLK(n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[14]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[15]  ( .D(n3765), 
        .CLK(n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[15]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[16]  ( .D(n3764), 
        .CLK(n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[16]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[17]  ( .D(n3763), 
        .CLK(n9177), .Q(CircularBuffer_sum_read_assign_reg_1610[17]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[18]  ( .D(n3762), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[18]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[19]  ( .D(n3761), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[19]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[20]  ( .D(n3760), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[20]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[21]  ( .D(n3759), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[21]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[22]  ( .D(n3758), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[22]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[23]  ( .D(n3757), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[23]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[24]  ( .D(n3756), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[24]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[25]  ( .D(n3755), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[25]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[26]  ( .D(n3754), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[26]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[27]  ( .D(n3753), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[27]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[28]  ( .D(n3752), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[28]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[29]  ( .D(n3751), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[29]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[30]  ( .D(n3750), 
        .CLK(n9176), .Q(CircularBuffer_sum_read_assign_reg_1610[30]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_reg_1610_reg[31]  ( .D(n3749), 
        .CLK(n9175), .Q(CircularBuffer_sum_read_assign_reg_1610[31]) );
  DFFPOSX1 \sum_reg_308_reg[0]  ( .D(n4471), .CLK(n9175), .Q(sum_reg_308[0])
         );
  DFFPOSX1 \recentVBools_sum_reg[0]  ( .D(n4439), .CLK(n9175), .Q(
        recentVBools_sum[0]) );
  DFFPOSX1 \sum_reg_308_reg[1]  ( .D(n4470), .CLK(n9175), .Q(sum_reg_308[1])
         );
  DFFPOSX1 \recentVBools_sum_reg[1]  ( .D(n4438), .CLK(n9175), .Q(
        recentVBools_sum[1]) );
  DFFPOSX1 \sum_reg_308_reg[2]  ( .D(n4469), .CLK(n9175), .Q(sum_reg_308[2])
         );
  DFFPOSX1 \recentVBools_sum_reg[2]  ( .D(n4437), .CLK(n9175), .Q(
        recentVBools_sum[2]) );
  DFFPOSX1 \sum_reg_308_reg[3]  ( .D(n4468), .CLK(n9175), .Q(sum_reg_308[3])
         );
  DFFPOSX1 \recentVBools_sum_reg[3]  ( .D(n4436), .CLK(n9175), .Q(
        recentVBools_sum[3]) );
  DFFPOSX1 \sum_reg_308_reg[4]  ( .D(n4467), .CLK(n9175), .Q(sum_reg_308[4])
         );
  DFFPOSX1 \recentVBools_sum_reg[4]  ( .D(n4435), .CLK(n9175), .Q(
        recentVBools_sum[4]) );
  DFFPOSX1 \sum_reg_308_reg[5]  ( .D(n4466), .CLK(n9175), .Q(sum_reg_308[5])
         );
  DFFPOSX1 \recentVBools_sum_reg[5]  ( .D(n4434), .CLK(n9175), .Q(
        recentVBools_sum[5]) );
  DFFPOSX1 \sum_reg_308_reg[6]  ( .D(n4465), .CLK(n9174), .Q(sum_reg_308[6])
         );
  DFFPOSX1 \recentVBools_sum_reg[6]  ( .D(n4433), .CLK(n9174), .Q(
        recentVBools_sum[6]) );
  DFFPOSX1 \sum_reg_308_reg[7]  ( .D(n4464), .CLK(n9174), .Q(sum_reg_308[7])
         );
  DFFPOSX1 \recentVBools_sum_reg[7]  ( .D(n4432), .CLK(n9174), .Q(
        recentVBools_sum[7]) );
  DFFPOSX1 \sum_reg_308_reg[8]  ( .D(n4463), .CLK(n9174), .Q(sum_reg_308[8])
         );
  DFFPOSX1 \recentVBools_sum_reg[8]  ( .D(n4431), .CLK(n9174), .Q(
        recentVBools_sum[8]) );
  DFFPOSX1 \sum_reg_308_reg[9]  ( .D(n4462), .CLK(n9174), .Q(sum_reg_308[9])
         );
  DFFPOSX1 \recentVBools_sum_reg[9]  ( .D(n4430), .CLK(n9174), .Q(
        recentVBools_sum[9]) );
  DFFPOSX1 \sum_reg_308_reg[10]  ( .D(n4461), .CLK(n9174), .Q(sum_reg_308[10])
         );
  DFFPOSX1 \recentVBools_sum_reg[10]  ( .D(n4429), .CLK(n9174), .Q(
        recentVBools_sum[10]) );
  DFFPOSX1 \sum_reg_308_reg[11]  ( .D(n4460), .CLK(n9174), .Q(sum_reg_308[11])
         );
  DFFPOSX1 \recentVBools_sum_reg[11]  ( .D(n4428), .CLK(n9174), .Q(
        recentVBools_sum[11]) );
  DFFPOSX1 \sum_reg_308_reg[12]  ( .D(n4459), .CLK(n9174), .Q(sum_reg_308[12])
         );
  DFFPOSX1 \recentVBools_sum_reg[12]  ( .D(n4427), .CLK(n9173), .Q(
        recentVBools_sum[12]) );
  DFFPOSX1 \sum_reg_308_reg[13]  ( .D(n4458), .CLK(n9173), .Q(sum_reg_308[13])
         );
  DFFPOSX1 \recentVBools_sum_reg[13]  ( .D(n4426), .CLK(n9173), .Q(
        recentVBools_sum[13]) );
  DFFPOSX1 \sum_reg_308_reg[14]  ( .D(n4457), .CLK(n9173), .Q(sum_reg_308[14])
         );
  DFFPOSX1 \recentVBools_sum_reg[14]  ( .D(n4425), .CLK(n9173), .Q(
        recentVBools_sum[14]) );
  DFFPOSX1 \sum_reg_308_reg[15]  ( .D(n4456), .CLK(n9173), .Q(sum_reg_308[15])
         );
  DFFPOSX1 \recentVBools_sum_reg[15]  ( .D(n4424), .CLK(n9173), .Q(
        recentVBools_sum[15]) );
  DFFPOSX1 \sum_reg_308_reg[16]  ( .D(n4455), .CLK(n9173), .Q(sum_reg_308[16])
         );
  DFFPOSX1 \recentVBools_sum_reg[16]  ( .D(n4423), .CLK(n9173), .Q(
        recentVBools_sum[16]) );
  DFFPOSX1 \sum_reg_308_reg[17]  ( .D(n4454), .CLK(n9173), .Q(sum_reg_308[17])
         );
  DFFPOSX1 \recentVBools_sum_reg[17]  ( .D(n4422), .CLK(n9173), .Q(
        recentVBools_sum[17]) );
  DFFPOSX1 \sum_reg_308_reg[18]  ( .D(n4453), .CLK(n9173), .Q(sum_reg_308[18])
         );
  DFFPOSX1 \recentVBools_sum_reg[18]  ( .D(n4421), .CLK(n9173), .Q(
        recentVBools_sum[18]) );
  DFFPOSX1 \sum_reg_308_reg[19]  ( .D(n4452), .CLK(n9172), .Q(sum_reg_308[19])
         );
  DFFPOSX1 \recentVBools_sum_reg[19]  ( .D(n4420), .CLK(n9172), .Q(
        recentVBools_sum[19]) );
  DFFPOSX1 \sum_reg_308_reg[20]  ( .D(n4451), .CLK(n9172), .Q(sum_reg_308[20])
         );
  DFFPOSX1 \recentVBools_sum_reg[20]  ( .D(n4419), .CLK(n9172), .Q(
        recentVBools_sum[20]) );
  DFFPOSX1 \sum_reg_308_reg[21]  ( .D(n4450), .CLK(n9172), .Q(sum_reg_308[21])
         );
  DFFPOSX1 \recentVBools_sum_reg[21]  ( .D(n4418), .CLK(n9172), .Q(
        recentVBools_sum[21]) );
  DFFPOSX1 \sum_reg_308_reg[22]  ( .D(n4449), .CLK(n9172), .Q(sum_reg_308[22])
         );
  DFFPOSX1 \recentVBools_sum_reg[22]  ( .D(n4417), .CLK(n9172), .Q(
        recentVBools_sum[22]) );
  DFFPOSX1 \sum_reg_308_reg[23]  ( .D(n4448), .CLK(n9172), .Q(sum_reg_308[23])
         );
  DFFPOSX1 \recentVBools_sum_reg[23]  ( .D(n4416), .CLK(n9172), .Q(
        recentVBools_sum[23]) );
  DFFPOSX1 \sum_reg_308_reg[24]  ( .D(n4447), .CLK(n9172), .Q(sum_reg_308[24])
         );
  DFFPOSX1 \recentVBools_sum_reg[24]  ( .D(n4415), .CLK(n9172), .Q(
        recentVBools_sum[24]) );
  DFFPOSX1 \sum_reg_308_reg[25]  ( .D(n4446), .CLK(n9172), .Q(sum_reg_308[25])
         );
  DFFPOSX1 \recentVBools_sum_reg[25]  ( .D(n4414), .CLK(n9171), .Q(
        recentVBools_sum[25]) );
  DFFPOSX1 \sum_reg_308_reg[26]  ( .D(n4445), .CLK(n9171), .Q(sum_reg_308[26])
         );
  DFFPOSX1 \recentVBools_sum_reg[26]  ( .D(n4413), .CLK(n9171), .Q(
        recentVBools_sum[26]) );
  DFFPOSX1 \sum_reg_308_reg[27]  ( .D(n4444), .CLK(n9171), .Q(sum_reg_308[27])
         );
  DFFPOSX1 \recentVBools_sum_reg[27]  ( .D(n4412), .CLK(n9171), .Q(
        recentVBools_sum[27]) );
  DFFPOSX1 \sum_reg_308_reg[28]  ( .D(n4443), .CLK(n9171), .Q(sum_reg_308[28])
         );
  DFFPOSX1 \recentVBools_sum_reg[28]  ( .D(n4411), .CLK(n9171), .Q(
        recentVBools_sum[28]) );
  DFFPOSX1 \sum_reg_308_reg[29]  ( .D(n4442), .CLK(n9171), .Q(sum_reg_308[29])
         );
  DFFPOSX1 \recentVBools_sum_reg[29]  ( .D(n4410), .CLK(n9171), .Q(
        recentVBools_sum[29]) );
  DFFPOSX1 \sum_reg_308_reg[30]  ( .D(n4441), .CLK(n9171), .Q(sum_reg_308[30])
         );
  DFFPOSX1 \recentVBools_sum_reg[30]  ( .D(n4409), .CLK(n9171), .Q(
        recentVBools_sum[30]) );
  DFFPOSX1 \sum_reg_308_reg[31]  ( .D(n4440), .CLK(n9171), .Q(sum_reg_308[31])
         );
  DFFPOSX1 \last_sample_is_V_V_loc_2_reg_358_reg[0]  ( .D(n4406), .CLK(n9171), 
        .Q(\last_sample_is_V_V_loc_2_reg_358[0] ) );
  DFFPOSX1 \last_sample_is_V_V_reg[0]  ( .D(n4407), .CLK(n9170), .Q(
        \last_sample_is_V_V[0] ) );
  DFFPOSX1 \recentVBools_sum_reg[31]  ( .D(n4408), .CLK(n9170), .Q(
        recentVBools_sum[31]) );
  DFFPOSX1 \ap_CS_fsm_reg[8]  ( .D(N106), .CLK(n9170), .Q(ap_CS_fsm[8]) );
  DFFPOSX1 \tmp_12_reg_1694_reg[0]  ( .D(n9471), .CLK(n9170), .Q(
        \tmp_12_reg_1694[0] ) );
  DFFPOSX1 \ap_CS_fsm_reg[9]  ( .D(N107), .CLK(n9170), .Q(ap_CS_fsm[9]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[30]  ( .D(n3747), 
        .CLK(n9170), .Q(CircularBuffer_sum_read_assign_1_reg_1705[30]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[29]  ( .D(n3746), 
        .CLK(n9170), .Q(CircularBuffer_sum_read_assign_1_reg_1705[29]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[28]  ( .D(n3745), 
        .CLK(n9170), .Q(CircularBuffer_sum_read_assign_1_reg_1705[28]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[27]  ( .D(n3744), 
        .CLK(n9170), .Q(CircularBuffer_sum_read_assign_1_reg_1705[27]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[26]  ( .D(n3743), 
        .CLK(n9170), .Q(CircularBuffer_sum_read_assign_1_reg_1705[26]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[25]  ( .D(n3742), 
        .CLK(n9170), .Q(CircularBuffer_sum_read_assign_1_reg_1705[25]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[24]  ( .D(n3741), 
        .CLK(n9170), .Q(CircularBuffer_sum_read_assign_1_reg_1705[24]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[23]  ( .D(n3740), 
        .CLK(n9170), .Q(CircularBuffer_sum_read_assign_1_reg_1705[23]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[22]  ( .D(n3739), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[22]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[21]  ( .D(n3738), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[21]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[20]  ( .D(n3737), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[20]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[19]  ( .D(n3736), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[19]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[18]  ( .D(n3735), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[18]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[17]  ( .D(n3734), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[17]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[16]  ( .D(n3733), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[16]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[15]  ( .D(n3732), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[15]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[14]  ( .D(n3731), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[14]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[13]  ( .D(n3730), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[13]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[12]  ( .D(n3729), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[12]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[11]  ( .D(n3728), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[11]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[10]  ( .D(n3727), 
        .CLK(n9169), .Q(CircularBuffer_sum_read_assign_1_reg_1705[10]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[9]  ( .D(n3726), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[9]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[8]  ( .D(n3725), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[8]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[7]  ( .D(n3724), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[7]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[6]  ( .D(n3723), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[6]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[5]  ( .D(n3722), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[5]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[4]  ( .D(n3721), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[4]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[3]  ( .D(n3720), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[3]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[2]  ( .D(n3719), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[2]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[1]  ( .D(n3718), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[1]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[0]  ( .D(n3717), 
        .CLK(n9168), .Q(CircularBuffer_sum_read_assign_1_reg_1705[0]) );
  DFFPOSX1 \recentABools_head_i_reg[0]  ( .D(n3716), .CLK(n9168), .Q(
        recentABools_head_i[0]) );
  DFFPOSX1 \recentABools_data_addr_reg_1689_reg[0]  ( .D(n3715), .CLK(n9168), 
        .Q(recentABools_data_addr_reg_1689[0]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[0]  ( .D(n3714), 
        .CLK(n9168), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[0]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[5]  ( .D(n3713), 
        .CLK(n9167), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[5]) );
  DFFPOSX1 \recentABools_head_i_reg[5]  ( .D(n3712), .CLK(n9167), .Q(
        recentABools_head_i[5]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[6]  ( .D(n3711), 
        .CLK(n9167), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[6]) );
  DFFPOSX1 \recentABools_head_i_reg[6]  ( .D(n3710), .CLK(n9167), .Q(
        recentABools_head_i[6]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[7]  ( .D(n3709), 
        .CLK(n9167), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[7]) );
  DFFPOSX1 \recentABools_head_i_reg[7]  ( .D(n3708), .CLK(n9167), .Q(
        recentABools_head_i[7]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[8]  ( .D(n3707), 
        .CLK(n9167), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[8]) );
  DFFPOSX1 \recentABools_head_i_reg[8]  ( .D(n3706), .CLK(n9167), .Q(
        recentABools_head_i[8]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[9]  ( .D(n3705), 
        .CLK(n9167), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[9]) );
  DFFPOSX1 \recentABools_head_i_reg[9]  ( .D(n3704), .CLK(n9167), .Q(
        recentABools_head_i[9]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[10]  ( .D(n3703), 
        .CLK(n9167), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[10]) );
  DFFPOSX1 \recentABools_head_i_reg[10]  ( .D(n3702), .CLK(n9167), .Q(
        recentABools_head_i[10]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[11]  ( .D(n3701), 
        .CLK(n9167), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[11]) );
  DFFPOSX1 \recentABools_head_i_reg[11]  ( .D(n3700), .CLK(n9166), .Q(
        recentABools_head_i[11]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[12]  ( .D(n3699), 
        .CLK(n9166), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[12]) );
  DFFPOSX1 \recentABools_head_i_reg[12]  ( .D(n3698), .CLK(n9166), .Q(
        recentABools_head_i[12]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[13]  ( .D(n3697), 
        .CLK(n9166), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[13]) );
  DFFPOSX1 \recentABools_head_i_reg[13]  ( .D(n3696), .CLK(n9166), .Q(
        recentABools_head_i[13]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[14]  ( .D(n3695), 
        .CLK(n9166), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[14]) );
  DFFPOSX1 \recentABools_head_i_reg[14]  ( .D(n3694), .CLK(n9166), .Q(
        recentABools_head_i[14]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[15]  ( .D(n3693), 
        .CLK(n9166), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[15]) );
  DFFPOSX1 \recentABools_head_i_reg[15]  ( .D(n3692), .CLK(n9166), .Q(
        recentABools_head_i[15]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[16]  ( .D(n3691), 
        .CLK(n9166), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[16]) );
  DFFPOSX1 \recentABools_head_i_reg[16]  ( .D(n3690), .CLK(n9166), .Q(
        recentABools_head_i[16]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[17]  ( .D(n3689), 
        .CLK(n9166), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[17]) );
  DFFPOSX1 \recentABools_head_i_reg[17]  ( .D(n3688), .CLK(n9166), .Q(
        recentABools_head_i[17]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[18]  ( .D(n3687), 
        .CLK(n9165), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[18]) );
  DFFPOSX1 \recentABools_head_i_reg[18]  ( .D(n3686), .CLK(n9165), .Q(
        recentABools_head_i[18]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[19]  ( .D(n3685), 
        .CLK(n9165), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[19]) );
  DFFPOSX1 \recentABools_head_i_reg[19]  ( .D(n3684), .CLK(n9165), .Q(
        recentABools_head_i[19]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[20]  ( .D(n3683), 
        .CLK(n9165), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[20]) );
  DFFPOSX1 \recentABools_head_i_reg[20]  ( .D(n3682), .CLK(n9165), .Q(
        recentABools_head_i[20]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[21]  ( .D(n3681), 
        .CLK(n9165), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[21]) );
  DFFPOSX1 \recentABools_head_i_reg[21]  ( .D(n3680), .CLK(n9165), .Q(
        recentABools_head_i[21]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[22]  ( .D(n3679), 
        .CLK(n9165), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[22]) );
  DFFPOSX1 \recentABools_head_i_reg[22]  ( .D(n3678), .CLK(n9165), .Q(
        recentABools_head_i[22]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[23]  ( .D(n3677), 
        .CLK(n9165), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[23]) );
  DFFPOSX1 \recentABools_head_i_reg[23]  ( .D(n3676), .CLK(n9165), .Q(
        recentABools_head_i[23]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[24]  ( .D(n3675), 
        .CLK(n9165), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[24]) );
  DFFPOSX1 \recentABools_head_i_reg[24]  ( .D(n3674), .CLK(n9164), .Q(
        recentABools_head_i[24]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[25]  ( .D(n3673), 
        .CLK(n9164), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[25]) );
  DFFPOSX1 \recentABools_head_i_reg[25]  ( .D(n3672), .CLK(n9164), .Q(
        recentABools_head_i[25]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[26]  ( .D(n3671), 
        .CLK(n9164), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[26]) );
  DFFPOSX1 \recentABools_head_i_reg[26]  ( .D(n3670), .CLK(n9164), .Q(
        recentABools_head_i[26]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[27]  ( .D(n3669), 
        .CLK(n9164), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[27]) );
  DFFPOSX1 \recentABools_head_i_reg[27]  ( .D(n3668), .CLK(n9164), .Q(
        recentABools_head_i[27]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[28]  ( .D(n3667), 
        .CLK(n9164), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[28]) );
  DFFPOSX1 \recentABools_head_i_reg[28]  ( .D(n3666), .CLK(n9164), .Q(
        recentABools_head_i[28]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[29]  ( .D(n3665), 
        .CLK(n9164), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[29]) );
  DFFPOSX1 \recentABools_head_i_reg[29]  ( .D(n3664), .CLK(n9164), .Q(
        recentABools_head_i[29]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[30]  ( .D(n3663), 
        .CLK(n9164), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[30]) );
  DFFPOSX1 \recentABools_head_i_reg[30]  ( .D(n3662), .CLK(n9164), .Q(
        recentABools_head_i[30]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[31]  ( .D(n3661), 
        .CLK(n9163), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[31]) );
  DFFPOSX1 \recentABools_head_i_reg[31]  ( .D(n3660), .CLK(n9163), .Q(
        recentABools_head_i[31]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[4]  ( .D(n7384), 
        .CLK(n9163), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[4]) );
  DFFPOSX1 \recentABools_head_i_reg[4]  ( .D(n3658), .CLK(n9163), .Q(
        recentABools_head_i[4]) );
  DFFPOSX1 \recentABools_data_addr_reg_1689_reg[4]  ( .D(n3657), .CLK(n9163), 
        .Q(recentABools_data_addr_reg_1689[4]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[3]  ( .D(n7565), 
        .CLK(n9163), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[3]) );
  DFFPOSX1 \recentABools_head_i_reg[3]  ( .D(n3655), .CLK(n9163), .Q(
        recentABools_head_i[3]) );
  DFFPOSX1 \recentABools_data_addr_reg_1689_reg[3]  ( .D(n3654), .CLK(n9163), 
        .Q(recentABools_data_addr_reg_1689[3]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[2]  ( .D(n7763), 
        .CLK(n9163), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[2]) );
  DFFPOSX1 \recentABools_head_i_reg[2]  ( .D(n3652), .CLK(n9163), .Q(
        recentABools_head_i[2]) );
  DFFPOSX1 \recentABools_data_addr_reg_1689_reg[2]  ( .D(n3651), .CLK(n9163), 
        .Q(recentABools_data_addr_reg_1689[2]) );
  DFFPOSX1 \CircularBuffer_head_i_read_ass_1_reg_1719_reg[1]  ( .D(n7981), 
        .CLK(n9163), .Q(CircularBuffer_head_i_read_ass_1_reg_1719[1]) );
  DFFPOSX1 \recentABools_head_i_reg[1]  ( .D(n3649), .CLK(n9163), .Q(
        recentABools_head_i[1]) );
  DFFPOSX1 \recentABools_data_addr_reg_1689_reg[1]  ( .D(n3648), .CLK(n9162), 
        .Q(recentABools_data_addr_reg_1689[1]) );
  DFFPOSX1 \VbeatFallDelay_reg[0]  ( .D(n3647), .CLK(n9162), .Q(
        VbeatFallDelay[0]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[0]  ( .D(n3646), .CLK(n9162), .Q(
        tmp_5_reg_1603[0]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[0]  ( .D(n4169), .CLK(n9162), .Q(
        VbeatFallDelay_new_1_reg_342[0]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[1]  ( .D(n3645), .CLK(n9162), .Q(
        tmp_5_reg_1603[1]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[1]  ( .D(n4170), .CLK(n9162), .Q(
        VbeatFallDelay_new_1_reg_342[1]) );
  DFFPOSX1 \VbeatFallDelay_reg[1]  ( .D(n3644), .CLK(n9162), .Q(
        VbeatFallDelay[1]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[2]  ( .D(n3643), .CLK(n9162), .Q(
        tmp_5_reg_1603[2]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[2]  ( .D(n4171), .CLK(n9162), .Q(
        VbeatFallDelay_new_1_reg_342[2]) );
  DFFPOSX1 \VbeatFallDelay_reg[2]  ( .D(n3642), .CLK(n9162), .Q(
        VbeatFallDelay[2]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[3]  ( .D(n3641), .CLK(n9162), .Q(
        tmp_5_reg_1603[3]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[3]  ( .D(n4172), .CLK(n9162), .Q(
        VbeatFallDelay_new_1_reg_342[3]) );
  DFFPOSX1 \VbeatFallDelay_reg[3]  ( .D(n3640), .CLK(n9162), .Q(
        VbeatFallDelay[3]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[4]  ( .D(n3639), .CLK(n9161), .Q(
        tmp_5_reg_1603[4]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[4]  ( .D(n4173), .CLK(n9161), .Q(
        VbeatFallDelay_new_1_reg_342[4]) );
  DFFPOSX1 \VbeatFallDelay_reg[4]  ( .D(n3638), .CLK(n9161), .Q(
        VbeatFallDelay[4]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[5]  ( .D(n3637), .CLK(n9161), .Q(
        tmp_5_reg_1603[5]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[5]  ( .D(n4174), .CLK(n9161), .Q(
        VbeatFallDelay_new_1_reg_342[5]) );
  DFFPOSX1 \VbeatFallDelay_reg[5]  ( .D(n3636), .CLK(n9161), .Q(
        VbeatFallDelay[5]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[6]  ( .D(n3635), .CLK(n9161), .Q(
        tmp_5_reg_1603[6]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[6]  ( .D(n4175), .CLK(n9161), .Q(
        VbeatFallDelay_new_1_reg_342[6]) );
  DFFPOSX1 \VbeatFallDelay_reg[6]  ( .D(n3634), .CLK(n9161), .Q(
        VbeatFallDelay[6]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[7]  ( .D(n3633), .CLK(n9161), .Q(
        tmp_5_reg_1603[7]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[7]  ( .D(n4176), .CLK(n9161), .Q(
        VbeatFallDelay_new_1_reg_342[7]) );
  DFFPOSX1 \VbeatFallDelay_reg[7]  ( .D(n3632), .CLK(n9161), .Q(
        VbeatFallDelay[7]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[8]  ( .D(n3631), .CLK(n9161), .Q(
        tmp_5_reg_1603[8]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[8]  ( .D(n4177), .CLK(n9160), .Q(
        VbeatFallDelay_new_1_reg_342[8]) );
  DFFPOSX1 \VbeatFallDelay_reg[8]  ( .D(n3630), .CLK(n9160), .Q(
        VbeatFallDelay[8]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[9]  ( .D(n3629), .CLK(n9160), .Q(
        tmp_5_reg_1603[9]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[9]  ( .D(n4178), .CLK(n9160), .Q(
        VbeatFallDelay_new_1_reg_342[9]) );
  DFFPOSX1 \VbeatFallDelay_reg[9]  ( .D(n3628), .CLK(n9160), .Q(
        VbeatFallDelay[9]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[10]  ( .D(n3627), .CLK(n9160), .Q(
        tmp_5_reg_1603[10]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[10]  ( .D(n4179), .CLK(n9160), 
        .Q(VbeatFallDelay_new_1_reg_342[10]) );
  DFFPOSX1 \VbeatFallDelay_reg[10]  ( .D(n3626), .CLK(n9160), .Q(
        VbeatFallDelay[10]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[11]  ( .D(n3625), .CLK(n9160), .Q(
        tmp_5_reg_1603[11]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[11]  ( .D(n4180), .CLK(n9160), 
        .Q(VbeatFallDelay_new_1_reg_342[11]) );
  DFFPOSX1 \VbeatFallDelay_reg[11]  ( .D(n3624), .CLK(n9160), .Q(
        VbeatFallDelay[11]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[12]  ( .D(n3623), .CLK(n9160), .Q(
        tmp_5_reg_1603[12]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[12]  ( .D(n4181), .CLK(n9160), 
        .Q(VbeatFallDelay_new_1_reg_342[12]) );
  DFFPOSX1 \VbeatFallDelay_reg[12]  ( .D(n3622), .CLK(n9159), .Q(
        VbeatFallDelay[12]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[13]  ( .D(n3621), .CLK(n9159), .Q(
        tmp_5_reg_1603[13]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[13]  ( .D(n4182), .CLK(n9159), 
        .Q(VbeatFallDelay_new_1_reg_342[13]) );
  DFFPOSX1 \VbeatFallDelay_reg[13]  ( .D(n3620), .CLK(n9159), .Q(
        VbeatFallDelay[13]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[14]  ( .D(n3619), .CLK(n9159), .Q(
        tmp_5_reg_1603[14]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[14]  ( .D(n4183), .CLK(n9159), 
        .Q(VbeatFallDelay_new_1_reg_342[14]) );
  DFFPOSX1 \VbeatFallDelay_reg[14]  ( .D(n3618), .CLK(n9159), .Q(
        VbeatFallDelay[14]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[15]  ( .D(n3617), .CLK(n9159), .Q(
        tmp_5_reg_1603[15]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[15]  ( .D(n4184), .CLK(n9159), 
        .Q(VbeatFallDelay_new_1_reg_342[15]) );
  DFFPOSX1 \VbeatFallDelay_reg[15]  ( .D(n3616), .CLK(n9159), .Q(
        VbeatFallDelay[15]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[16]  ( .D(n3615), .CLK(n9159), .Q(
        tmp_5_reg_1603[16]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[16]  ( .D(n4185), .CLK(n9159), 
        .Q(VbeatFallDelay_new_1_reg_342[16]) );
  DFFPOSX1 \VbeatFallDelay_reg[16]  ( .D(n3614), .CLK(n9159), .Q(
        VbeatFallDelay[16]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[17]  ( .D(n3613), .CLK(n9158), .Q(
        tmp_5_reg_1603[17]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[17]  ( .D(n4186), .CLK(n9158), 
        .Q(VbeatFallDelay_new_1_reg_342[17]) );
  DFFPOSX1 \VbeatFallDelay_reg[17]  ( .D(n3612), .CLK(n9158), .Q(
        VbeatFallDelay[17]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[18]  ( .D(n3611), .CLK(n9158), .Q(
        tmp_5_reg_1603[18]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[18]  ( .D(n4187), .CLK(n9158), 
        .Q(VbeatFallDelay_new_1_reg_342[18]) );
  DFFPOSX1 \VbeatFallDelay_reg[18]  ( .D(n3610), .CLK(n9158), .Q(
        VbeatFallDelay[18]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[19]  ( .D(n3609), .CLK(n9158), .Q(
        tmp_5_reg_1603[19]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[19]  ( .D(n4188), .CLK(n9158), 
        .Q(VbeatFallDelay_new_1_reg_342[19]) );
  DFFPOSX1 \VbeatFallDelay_reg[19]  ( .D(n3608), .CLK(n9158), .Q(
        VbeatFallDelay[19]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[20]  ( .D(n3607), .CLK(n9158), .Q(
        tmp_5_reg_1603[20]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[20]  ( .D(n4189), .CLK(n9158), 
        .Q(VbeatFallDelay_new_1_reg_342[20]) );
  DFFPOSX1 \VbeatFallDelay_reg[20]  ( .D(n3606), .CLK(n9158), .Q(
        VbeatFallDelay[20]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[21]  ( .D(n3605), .CLK(n9158), .Q(
        tmp_5_reg_1603[21]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[21]  ( .D(n4190), .CLK(n9157), 
        .Q(VbeatFallDelay_new_1_reg_342[21]) );
  DFFPOSX1 \VbeatFallDelay_reg[21]  ( .D(n3604), .CLK(n9157), .Q(
        VbeatFallDelay[21]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[22]  ( .D(n3603), .CLK(n9157), .Q(
        tmp_5_reg_1603[22]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[22]  ( .D(n4191), .CLK(n9157), 
        .Q(VbeatFallDelay_new_1_reg_342[22]) );
  DFFPOSX1 \VbeatFallDelay_reg[22]  ( .D(n3602), .CLK(n9157), .Q(
        VbeatFallDelay[22]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[23]  ( .D(n3601), .CLK(n9157), .Q(
        tmp_5_reg_1603[23]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[23]  ( .D(n4192), .CLK(n9157), 
        .Q(VbeatFallDelay_new_1_reg_342[23]) );
  DFFPOSX1 \VbeatFallDelay_reg[23]  ( .D(n3600), .CLK(n9157), .Q(
        VbeatFallDelay[23]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[24]  ( .D(n3599), .CLK(n9157), .Q(
        tmp_5_reg_1603[24]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[24]  ( .D(n4193), .CLK(n9157), 
        .Q(VbeatFallDelay_new_1_reg_342[24]) );
  DFFPOSX1 \VbeatFallDelay_reg[24]  ( .D(n3598), .CLK(n9157), .Q(
        VbeatFallDelay[24]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[25]  ( .D(n3597), .CLK(n9157), .Q(
        tmp_5_reg_1603[25]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[25]  ( .D(n4194), .CLK(n9157), 
        .Q(VbeatFallDelay_new_1_reg_342[25]) );
  DFFPOSX1 \VbeatFallDelay_reg[25]  ( .D(n3596), .CLK(n9156), .Q(
        VbeatFallDelay[25]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[26]  ( .D(n3595), .CLK(n9156), .Q(
        tmp_5_reg_1603[26]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[26]  ( .D(n4195), .CLK(n9156), 
        .Q(VbeatFallDelay_new_1_reg_342[26]) );
  DFFPOSX1 \VbeatFallDelay_reg[26]  ( .D(n3594), .CLK(n9156), .Q(
        VbeatFallDelay[26]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[27]  ( .D(n3593), .CLK(n9156), .Q(
        tmp_5_reg_1603[27]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[27]  ( .D(n4196), .CLK(n9156), 
        .Q(VbeatFallDelay_new_1_reg_342[27]) );
  DFFPOSX1 \VbeatFallDelay_reg[27]  ( .D(n3592), .CLK(n9156), .Q(
        VbeatFallDelay[27]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[28]  ( .D(n3591), .CLK(n9156), .Q(
        tmp_5_reg_1603[28]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[28]  ( .D(n4197), .CLK(n9156), 
        .Q(VbeatFallDelay_new_1_reg_342[28]) );
  DFFPOSX1 \VbeatFallDelay_reg[28]  ( .D(n3590), .CLK(n9156), .Q(
        VbeatFallDelay[28]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[29]  ( .D(n3589), .CLK(n9156), .Q(
        tmp_5_reg_1603[29]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[29]  ( .D(n4198), .CLK(n9156), 
        .Q(VbeatFallDelay_new_1_reg_342[29]) );
  DFFPOSX1 \VbeatFallDelay_reg[29]  ( .D(n3588), .CLK(n9156), .Q(
        VbeatFallDelay[29]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[30]  ( .D(n3587), .CLK(n9155), .Q(
        tmp_5_reg_1603[30]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[30]  ( .D(n4199), .CLK(n9155), 
        .Q(VbeatFallDelay_new_1_reg_342[30]) );
  DFFPOSX1 \VbeatFallDelay_reg[30]  ( .D(n3586), .CLK(n9155), .Q(
        VbeatFallDelay[30]) );
  DFFPOSX1 \tmp_5_reg_1603_reg[31]  ( .D(n3585), .CLK(n9155), .Q(
        tmp_5_reg_1603[31]) );
  DFFPOSX1 \VbeatFallDelay_new_1_reg_342_reg[31]  ( .D(n4200), .CLK(n9155), 
        .Q(VbeatFallDelay_new_1_reg_342[31]) );
  DFFPOSX1 \VbeatFallDelay_reg[31]  ( .D(n3584), .CLK(n9155), .Q(
        VbeatFallDelay[31]) );
  DFFPOSX1 \VbeatDelay_reg[3]  ( .D(n3583), .CLK(n9155), .Q(VbeatDelay[3]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[0]  ( .D(n3582), .CLK(n9155), .Q(
        tmp_4_reg_1596[0]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[0]  ( .D(n4405), .CLK(n9155), .Q(
        VbeatDelay_new_1_reg_326[0]) );
  DFFPOSX1 \VbeatDelay_reg[0]  ( .D(n3581), .CLK(n9155), .Q(VbeatDelay[0]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[1]  ( .D(n3580), .CLK(n9155), .Q(
        tmp_4_reg_1596[1]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[1]  ( .D(n4404), .CLK(n9155), .Q(
        VbeatDelay_new_1_reg_326[1]) );
  DFFPOSX1 \VbeatDelay_reg[1]  ( .D(n3579), .CLK(n9155), .Q(VbeatDelay[1]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[2]  ( .D(n3578), .CLK(n9154), .Q(
        tmp_4_reg_1596[2]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[2]  ( .D(n4403), .CLK(n9154), .Q(
        VbeatDelay_new_1_reg_326[2]) );
  DFFPOSX1 \VbeatDelay_reg[2]  ( .D(n3577), .CLK(n9154), .Q(VbeatDelay[2]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[3]  ( .D(n3576), .CLK(n9154), .Q(
        tmp_4_reg_1596[3]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[3]  ( .D(n4402), .CLK(n9154), .Q(
        VbeatDelay_new_1_reg_326[3]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[4]  ( .D(n3575), .CLK(n9154), .Q(
        tmp_4_reg_1596[4]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[4]  ( .D(n4401), .CLK(n9154), .Q(
        VbeatDelay_new_1_reg_326[4]) );
  DFFPOSX1 \VbeatDelay_reg[4]  ( .D(n3574), .CLK(n9154), .Q(VbeatDelay[4]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[5]  ( .D(n3573), .CLK(n9154), .Q(
        tmp_4_reg_1596[5]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[5]  ( .D(n4400), .CLK(n9154), .Q(
        VbeatDelay_new_1_reg_326[5]) );
  DFFPOSX1 \VbeatDelay_reg[5]  ( .D(n3572), .CLK(n9154), .Q(VbeatDelay[5]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[6]  ( .D(n3571), .CLK(n9154), .Q(
        tmp_4_reg_1596[6]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[6]  ( .D(n4399), .CLK(n9154), .Q(
        VbeatDelay_new_1_reg_326[6]) );
  DFFPOSX1 \VbeatDelay_reg[6]  ( .D(n3570), .CLK(n9153), .Q(VbeatDelay[6]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[7]  ( .D(n3569), .CLK(n9153), .Q(
        tmp_4_reg_1596[7]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[7]  ( .D(n4398), .CLK(n9153), .Q(
        VbeatDelay_new_1_reg_326[7]) );
  DFFPOSX1 \VbeatDelay_reg[7]  ( .D(n3568), .CLK(n9153), .Q(VbeatDelay[7]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[8]  ( .D(n3567), .CLK(n9153), .Q(
        tmp_4_reg_1596[8]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[8]  ( .D(n4397), .CLK(n9153), .Q(
        VbeatDelay_new_1_reg_326[8]) );
  DFFPOSX1 \VbeatDelay_reg[8]  ( .D(n3566), .CLK(n9153), .Q(VbeatDelay[8]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[9]  ( .D(n3565), .CLK(n9153), .Q(
        tmp_4_reg_1596[9]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[9]  ( .D(n4396), .CLK(n9153), .Q(
        VbeatDelay_new_1_reg_326[9]) );
  DFFPOSX1 \VbeatDelay_reg[9]  ( .D(n3564), .CLK(n9153), .Q(VbeatDelay[9]) );
  DFFPOSX1 \tmp_4_reg_1596_reg[10]  ( .D(n3563), .CLK(n9153), .Q(
        tmp_4_reg_1596[10]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[10]  ( .D(n4395), .CLK(n9153), .Q(
        VbeatDelay_new_1_reg_326[10]) );
  DFFPOSX1 \VbeatDelay_reg[10]  ( .D(n3562), .CLK(n9153), .Q(VbeatDelay[10])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[11]  ( .D(n3561), .CLK(n9152), .Q(
        tmp_4_reg_1596[11]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[11]  ( .D(n4394), .CLK(n9152), .Q(
        VbeatDelay_new_1_reg_326[11]) );
  DFFPOSX1 \VbeatDelay_reg[11]  ( .D(n3560), .CLK(n9152), .Q(VbeatDelay[11])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[12]  ( .D(n3559), .CLK(n9152), .Q(
        tmp_4_reg_1596[12]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[12]  ( .D(n4393), .CLK(n9152), .Q(
        VbeatDelay_new_1_reg_326[12]) );
  DFFPOSX1 \VbeatDelay_reg[12]  ( .D(n3558), .CLK(n9152), .Q(VbeatDelay[12])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[13]  ( .D(n3557), .CLK(n9152), .Q(
        tmp_4_reg_1596[13]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[13]  ( .D(n4392), .CLK(n9152), .Q(
        VbeatDelay_new_1_reg_326[13]) );
  DFFPOSX1 \VbeatDelay_reg[13]  ( .D(n3556), .CLK(n9152), .Q(VbeatDelay[13])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[14]  ( .D(n3555), .CLK(n9152), .Q(
        tmp_4_reg_1596[14]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[14]  ( .D(n4391), .CLK(n9152), .Q(
        VbeatDelay_new_1_reg_326[14]) );
  DFFPOSX1 \VbeatDelay_reg[14]  ( .D(n3554), .CLK(n9152), .Q(VbeatDelay[14])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[15]  ( .D(n3553), .CLK(n9152), .Q(
        tmp_4_reg_1596[15]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[15]  ( .D(n4390), .CLK(n9151), .Q(
        VbeatDelay_new_1_reg_326[15]) );
  DFFPOSX1 \VbeatDelay_reg[15]  ( .D(n3552), .CLK(n9151), .Q(VbeatDelay[15])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[16]  ( .D(n3551), .CLK(n9151), .Q(
        tmp_4_reg_1596[16]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[16]  ( .D(n4389), .CLK(n9151), .Q(
        VbeatDelay_new_1_reg_326[16]) );
  DFFPOSX1 \VbeatDelay_reg[16]  ( .D(n3550), .CLK(n9151), .Q(VbeatDelay[16])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[17]  ( .D(n3549), .CLK(n9151), .Q(
        tmp_4_reg_1596[17]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[17]  ( .D(n4388), .CLK(n9151), .Q(
        VbeatDelay_new_1_reg_326[17]) );
  DFFPOSX1 \VbeatDelay_reg[17]  ( .D(n3548), .CLK(n9151), .Q(VbeatDelay[17])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[18]  ( .D(n3547), .CLK(n9151), .Q(
        tmp_4_reg_1596[18]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[18]  ( .D(n4387), .CLK(n9151), .Q(
        VbeatDelay_new_1_reg_326[18]) );
  DFFPOSX1 \VbeatDelay_reg[18]  ( .D(n3546), .CLK(n9151), .Q(VbeatDelay[18])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[19]  ( .D(n3545), .CLK(n9151), .Q(
        tmp_4_reg_1596[19]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[19]  ( .D(n4386), .CLK(n9151), .Q(
        VbeatDelay_new_1_reg_326[19]) );
  DFFPOSX1 \VbeatDelay_reg[19]  ( .D(n3544), .CLK(n9150), .Q(VbeatDelay[19])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[20]  ( .D(n3543), .CLK(n9150), .Q(
        tmp_4_reg_1596[20]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[20]  ( .D(n4385), .CLK(n9150), .Q(
        VbeatDelay_new_1_reg_326[20]) );
  DFFPOSX1 \VbeatDelay_reg[20]  ( .D(n3542), .CLK(n9150), .Q(VbeatDelay[20])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[21]  ( .D(n3541), .CLK(n9150), .Q(
        tmp_4_reg_1596[21]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[21]  ( .D(n4384), .CLK(n9150), .Q(
        VbeatDelay_new_1_reg_326[21]) );
  DFFPOSX1 \VbeatDelay_reg[21]  ( .D(n3540), .CLK(n9150), .Q(VbeatDelay[21])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[22]  ( .D(n3539), .CLK(n9150), .Q(
        tmp_4_reg_1596[22]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[22]  ( .D(n4383), .CLK(n9150), .Q(
        VbeatDelay_new_1_reg_326[22]) );
  DFFPOSX1 \VbeatDelay_reg[22]  ( .D(n3538), .CLK(n9150), .Q(VbeatDelay[22])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[23]  ( .D(n3537), .CLK(n9150), .Q(
        tmp_4_reg_1596[23]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[23]  ( .D(n4382), .CLK(n9150), .Q(
        VbeatDelay_new_1_reg_326[23]) );
  DFFPOSX1 \VbeatDelay_reg[23]  ( .D(n3536), .CLK(n9150), .Q(VbeatDelay[23])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[24]  ( .D(n3535), .CLK(n9149), .Q(
        tmp_4_reg_1596[24]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[24]  ( .D(n4381), .CLK(n9149), .Q(
        VbeatDelay_new_1_reg_326[24]) );
  DFFPOSX1 \VbeatDelay_reg[24]  ( .D(n3534), .CLK(n9149), .Q(VbeatDelay[24])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[25]  ( .D(n3533), .CLK(n9149), .Q(
        tmp_4_reg_1596[25]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[25]  ( .D(n4380), .CLK(n9149), .Q(
        VbeatDelay_new_1_reg_326[25]) );
  DFFPOSX1 \VbeatDelay_reg[25]  ( .D(n3532), .CLK(n9149), .Q(VbeatDelay[25])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[26]  ( .D(n3531), .CLK(n9149), .Q(
        tmp_4_reg_1596[26]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[26]  ( .D(n4379), .CLK(n9149), .Q(
        VbeatDelay_new_1_reg_326[26]) );
  DFFPOSX1 \VbeatDelay_reg[26]  ( .D(n3530), .CLK(n9149), .Q(VbeatDelay[26])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[27]  ( .D(n3529), .CLK(n9149), .Q(
        tmp_4_reg_1596[27]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[27]  ( .D(n4378), .CLK(n9149), .Q(
        VbeatDelay_new_1_reg_326[27]) );
  DFFPOSX1 \VbeatDelay_reg[27]  ( .D(n3528), .CLK(n9149), .Q(VbeatDelay[27])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[28]  ( .D(n3527), .CLK(n9149), .Q(
        tmp_4_reg_1596[28]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[28]  ( .D(n4377), .CLK(n9148), .Q(
        VbeatDelay_new_1_reg_326[28]) );
  DFFPOSX1 \VbeatDelay_reg[28]  ( .D(n3526), .CLK(n9148), .Q(VbeatDelay[28])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[29]  ( .D(n3525), .CLK(n9148), .Q(
        tmp_4_reg_1596[29]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[29]  ( .D(n4376), .CLK(n9148), .Q(
        VbeatDelay_new_1_reg_326[29]) );
  DFFPOSX1 \VbeatDelay_reg[29]  ( .D(n3524), .CLK(n9148), .Q(VbeatDelay[29])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[30]  ( .D(n3523), .CLK(n9148), .Q(
        tmp_4_reg_1596[30]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[30]  ( .D(n4375), .CLK(n9148), .Q(
        VbeatDelay_new_1_reg_326[30]) );
  DFFPOSX1 \VbeatDelay_reg[30]  ( .D(n3522), .CLK(n9148), .Q(VbeatDelay[30])
         );
  DFFPOSX1 \tmp_4_reg_1596_reg[31]  ( .D(n3521), .CLK(n9148), .Q(
        tmp_4_reg_1596[31]) );
  DFFPOSX1 \VbeatDelay_new_1_reg_326_reg[31]  ( .D(n4374), .CLK(n9148), .Q(
        VbeatDelay_new_1_reg_326[31]) );
  DFFPOSX1 \VbeatDelay_reg[31]  ( .D(n3520), .CLK(n9148), .Q(VbeatDelay[31])
         );
  DFFPOSX1 \ap_CS_fsm_reg[10]  ( .D(N108), .CLK(n9148), .Q(ap_CS_fsm[10]) );
  DFFPOSX1 \ap_CS_fsm_reg[11]  ( .D(N109), .CLK(n9148), .Q(ap_CS_fsm[11]) );
  DFFPOSX1 \ap_CS_fsm_reg[12]  ( .D(n4760), .CLK(n9147), .Q(ap_CS_fsm[12]) );
  DFFPOSX1 \recentABools_len_reg[0]  ( .D(n4340), .CLK(n9147), .Q(
        recentABools_len[0]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[0]  ( .D(n3519), 
        .CLK(n9147), .Q(CircularBuffer_len_write_assig_3_fu_1249_p2[0]) );
  DFFPOSX1 \tmp_13_reg_1725_reg[0]  ( .D(n3518), .CLK(n9147), .Q(
        \tmp_13_reg_1725[0] ) );
  DFFPOSX1 \sum_1_reg_376_reg[0]  ( .D(n4308), .CLK(n9147), .Q(
        sum_1_reg_376[0]) );
  DFFPOSX1 \recentABools_sum_reg[0]  ( .D(n4342), .CLK(n9147), .Q(
        recentABools_sum[0]) );
  DFFPOSX1 \sum_1_reg_376_reg[1]  ( .D(n4307), .CLK(n9147), .Q(
        sum_1_reg_376[1]) );
  DFFPOSX1 \recentABools_sum_reg[1]  ( .D(n4343), .CLK(n9147), .Q(
        recentABools_sum[1]) );
  DFFPOSX1 \sum_1_reg_376_reg[2]  ( .D(n4306), .CLK(n9147), .Q(
        sum_1_reg_376[2]) );
  DFFPOSX1 \recentABools_sum_reg[2]  ( .D(n4344), .CLK(n9147), .Q(
        recentABools_sum[2]) );
  DFFPOSX1 \sum_1_reg_376_reg[3]  ( .D(n4305), .CLK(n9147), .Q(
        sum_1_reg_376[3]) );
  DFFPOSX1 \recentABools_sum_reg[3]  ( .D(n4345), .CLK(n9147), .Q(
        recentABools_sum[3]) );
  DFFPOSX1 \sum_1_reg_376_reg[4]  ( .D(n4304), .CLK(n9147), .Q(
        sum_1_reg_376[4]) );
  DFFPOSX1 \recentABools_sum_reg[4]  ( .D(n4346), .CLK(n9146), .Q(
        recentABools_sum[4]) );
  DFFPOSX1 \sum_1_reg_376_reg[5]  ( .D(n4303), .CLK(n9146), .Q(
        sum_1_reg_376[5]) );
  DFFPOSX1 \recentABools_sum_reg[5]  ( .D(n4347), .CLK(n9146), .Q(
        recentABools_sum[5]) );
  DFFPOSX1 \sum_1_reg_376_reg[6]  ( .D(n4302), .CLK(n9146), .Q(
        sum_1_reg_376[6]) );
  DFFPOSX1 \recentABools_sum_reg[6]  ( .D(n4348), .CLK(n9146), .Q(
        recentABools_sum[6]) );
  DFFPOSX1 \sum_1_reg_376_reg[7]  ( .D(n4301), .CLK(n9146), .Q(
        sum_1_reg_376[7]) );
  DFFPOSX1 \recentABools_sum_reg[7]  ( .D(n4349), .CLK(n9146), .Q(
        recentABools_sum[7]) );
  DFFPOSX1 \sum_1_reg_376_reg[8]  ( .D(n4300), .CLK(n9146), .Q(
        sum_1_reg_376[8]) );
  DFFPOSX1 \recentABools_sum_reg[8]  ( .D(n4350), .CLK(n9146), .Q(
        recentABools_sum[8]) );
  DFFPOSX1 \sum_1_reg_376_reg[9]  ( .D(n4299), .CLK(n9146), .Q(
        sum_1_reg_376[9]) );
  DFFPOSX1 \recentABools_sum_reg[9]  ( .D(n4351), .CLK(n9146), .Q(
        recentABools_sum[9]) );
  DFFPOSX1 \sum_1_reg_376_reg[10]  ( .D(n4298), .CLK(n9146), .Q(
        sum_1_reg_376[10]) );
  DFFPOSX1 \recentABools_sum_reg[10]  ( .D(n4352), .CLK(n9146), .Q(
        recentABools_sum[10]) );
  DFFPOSX1 \sum_1_reg_376_reg[11]  ( .D(n4297), .CLK(n9145), .Q(
        sum_1_reg_376[11]) );
  DFFPOSX1 \recentABools_sum_reg[11]  ( .D(n4353), .CLK(n9145), .Q(
        recentABools_sum[11]) );
  DFFPOSX1 \sum_1_reg_376_reg[12]  ( .D(n4296), .CLK(n9145), .Q(
        sum_1_reg_376[12]) );
  DFFPOSX1 \recentABools_sum_reg[12]  ( .D(n4354), .CLK(n9145), .Q(
        recentABools_sum[12]) );
  DFFPOSX1 \sum_1_reg_376_reg[13]  ( .D(n4295), .CLK(n9145), .Q(
        sum_1_reg_376[13]) );
  DFFPOSX1 \recentABools_sum_reg[13]  ( .D(n4355), .CLK(n9145), .Q(
        recentABools_sum[13]) );
  DFFPOSX1 \sum_1_reg_376_reg[14]  ( .D(n4294), .CLK(n9145), .Q(
        sum_1_reg_376[14]) );
  DFFPOSX1 \recentABools_sum_reg[14]  ( .D(n4356), .CLK(n9145), .Q(
        recentABools_sum[14]) );
  DFFPOSX1 \sum_1_reg_376_reg[15]  ( .D(n4293), .CLK(n9145), .Q(
        sum_1_reg_376[15]) );
  DFFPOSX1 \recentABools_sum_reg[15]  ( .D(n4357), .CLK(n9145), .Q(
        recentABools_sum[15]) );
  DFFPOSX1 \sum_1_reg_376_reg[16]  ( .D(n4292), .CLK(n9145), .Q(
        sum_1_reg_376[16]) );
  DFFPOSX1 \recentABools_sum_reg[16]  ( .D(n4358), .CLK(n9145), .Q(
        recentABools_sum[16]) );
  DFFPOSX1 \sum_1_reg_376_reg[17]  ( .D(n4291), .CLK(n9145), .Q(
        sum_1_reg_376[17]) );
  DFFPOSX1 \recentABools_sum_reg[17]  ( .D(n4359), .CLK(n9144), .Q(
        recentABools_sum[17]) );
  DFFPOSX1 \sum_1_reg_376_reg[18]  ( .D(n4290), .CLK(n9144), .Q(
        sum_1_reg_376[18]) );
  DFFPOSX1 \recentABools_sum_reg[18]  ( .D(n4360), .CLK(n9144), .Q(
        recentABools_sum[18]) );
  DFFPOSX1 \sum_1_reg_376_reg[19]  ( .D(n4289), .CLK(n9144), .Q(
        sum_1_reg_376[19]) );
  DFFPOSX1 \recentABools_sum_reg[19]  ( .D(n4361), .CLK(n9144), .Q(
        recentABools_sum[19]) );
  DFFPOSX1 \sum_1_reg_376_reg[20]  ( .D(n4288), .CLK(n9144), .Q(
        sum_1_reg_376[20]) );
  DFFPOSX1 \recentABools_sum_reg[20]  ( .D(n4362), .CLK(n9144), .Q(
        recentABools_sum[20]) );
  DFFPOSX1 \sum_1_reg_376_reg[21]  ( .D(n4287), .CLK(n9144), .Q(
        sum_1_reg_376[21]) );
  DFFPOSX1 \recentABools_sum_reg[21]  ( .D(n4363), .CLK(n9144), .Q(
        recentABools_sum[21]) );
  DFFPOSX1 \sum_1_reg_376_reg[22]  ( .D(n4286), .CLK(n9144), .Q(
        sum_1_reg_376[22]) );
  DFFPOSX1 \recentABools_sum_reg[22]  ( .D(n4364), .CLK(n9144), .Q(
        recentABools_sum[22]) );
  DFFPOSX1 \sum_1_reg_376_reg[23]  ( .D(n4285), .CLK(n9144), .Q(
        sum_1_reg_376[23]) );
  DFFPOSX1 \recentABools_sum_reg[23]  ( .D(n4365), .CLK(n9144), .Q(
        recentABools_sum[23]) );
  DFFPOSX1 \sum_1_reg_376_reg[24]  ( .D(n4284), .CLK(n9143), .Q(
        sum_1_reg_376[24]) );
  DFFPOSX1 \recentABools_sum_reg[24]  ( .D(n4366), .CLK(n9143), .Q(
        recentABools_sum[24]) );
  DFFPOSX1 \sum_1_reg_376_reg[25]  ( .D(n4283), .CLK(n9143), .Q(
        sum_1_reg_376[25]) );
  DFFPOSX1 \recentABools_sum_reg[25]  ( .D(n4367), .CLK(n9143), .Q(
        recentABools_sum[25]) );
  DFFPOSX1 \sum_1_reg_376_reg[26]  ( .D(n4282), .CLK(n9143), .Q(
        sum_1_reg_376[26]) );
  DFFPOSX1 \recentABools_sum_reg[26]  ( .D(n4368), .CLK(n9143), .Q(
        recentABools_sum[26]) );
  DFFPOSX1 \sum_1_reg_376_reg[27]  ( .D(n4281), .CLK(n9143), .Q(
        sum_1_reg_376[27]) );
  DFFPOSX1 \recentABools_sum_reg[27]  ( .D(n4369), .CLK(n9143), .Q(
        recentABools_sum[27]) );
  DFFPOSX1 \sum_1_reg_376_reg[28]  ( .D(n4280), .CLK(n9143), .Q(
        sum_1_reg_376[28]) );
  DFFPOSX1 \recentABools_sum_reg[28]  ( .D(n4370), .CLK(n9143), .Q(
        recentABools_sum[28]) );
  DFFPOSX1 \sum_1_reg_376_reg[29]  ( .D(n4279), .CLK(n9143), .Q(
        sum_1_reg_376[29]) );
  DFFPOSX1 \recentABools_sum_reg[29]  ( .D(n4371), .CLK(n9143), .Q(
        recentABools_sum[29]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[30]  ( .D(n4246), .CLK(n9143), 
        .Q(recentABools_len_new_reg_385[30]) );
  DFFPOSX1 \recentABools_len_reg[30]  ( .D(n4310), .CLK(n9142), .Q(
        recentABools_len[30]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[1]  ( .D(n3517), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[1]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[2]  ( .D(n3516), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[2]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[3]  ( .D(n3515), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[3]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[4]  ( .D(n3514), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[4]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[5]  ( .D(n3513), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[5]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[6]  ( .D(n3512), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[6]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[7]  ( .D(n3511), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[7]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[8]  ( .D(n3510), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[8]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[9]  ( .D(n3509), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[9]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[10]  ( .D(n3508), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[10]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[11]  ( .D(n3507), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[11]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[12]  ( .D(n3506), 
        .CLK(n9142), .Q(CircularBuffer_len_read_assign_3_reg_1711[12]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[13]  ( .D(n3505), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[13]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[14]  ( .D(n3504), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[14]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[15]  ( .D(n3503), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[15]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[16]  ( .D(n3502), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[16]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[17]  ( .D(n3501), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[17]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[18]  ( .D(n3500), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[18]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[19]  ( .D(n3499), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[19]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[20]  ( .D(n3498), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[20]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[21]  ( .D(n3497), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[21]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[22]  ( .D(n3496), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[22]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[23]  ( .D(n3495), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[23]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[24]  ( .D(n3494), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[24]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[25]  ( .D(n3493), 
        .CLK(n9141), .Q(CircularBuffer_len_read_assign_3_reg_1711[25]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[26]  ( .D(n3492), 
        .CLK(n9140), .Q(CircularBuffer_len_read_assign_3_reg_1711[26]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[27]  ( .D(n3491), 
        .CLK(n9140), .Q(CircularBuffer_len_read_assign_3_reg_1711[27]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[28]  ( .D(n3490), 
        .CLK(n9140), .Q(CircularBuffer_len_read_assign_3_reg_1711[28]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[29]  ( .D(n3489), 
        .CLK(n9140), .Q(CircularBuffer_len_read_assign_3_reg_1711[29]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[30]  ( .D(n3488), 
        .CLK(n9140), .Q(CircularBuffer_len_read_assign_3_reg_1711[30]) );
  DFFPOSX1 \CircularBuffer_len_read_assign_3_reg_1711_reg[31]  ( .D(n3487), 
        .CLK(n9140), .Q(CircularBuffer_len_read_assign_3_reg_1711[31]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[1]  ( .D(n4275), .CLK(n9140), .Q(
        recentABools_len_new_reg_385[1]) );
  DFFPOSX1 \recentABools_len_reg[1]  ( .D(n4339), .CLK(n9140), .Q(
        recentABools_len[1]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[2]  ( .D(n4274), .CLK(n9140), .Q(
        recentABools_len_new_reg_385[2]) );
  DFFPOSX1 \recentABools_len_reg[2]  ( .D(n4338), .CLK(n9140), .Q(
        recentABools_len[2]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[3]  ( .D(n4273), .CLK(n9140), .Q(
        recentABools_len_new_reg_385[3]) );
  DFFPOSX1 \recentABools_len_reg[3]  ( .D(n4337), .CLK(n9140), .Q(
        recentABools_len[3]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[4]  ( .D(n4272), .CLK(n9140), .Q(
        recentABools_len_new_reg_385[4]) );
  DFFPOSX1 \recentABools_len_reg[4]  ( .D(n4336), .CLK(n9139), .Q(
        recentABools_len[4]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[5]  ( .D(n4271), .CLK(n9139), .Q(
        recentABools_len_new_reg_385[5]) );
  DFFPOSX1 \recentABools_len_reg[5]  ( .D(n4335), .CLK(n9139), .Q(
        recentABools_len[5]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[6]  ( .D(n4270), .CLK(n9139), .Q(
        recentABools_len_new_reg_385[6]) );
  DFFPOSX1 \recentABools_len_reg[6]  ( .D(n4334), .CLK(n9139), .Q(
        recentABools_len[6]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[7]  ( .D(n4269), .CLK(n9139), .Q(
        recentABools_len_new_reg_385[7]) );
  DFFPOSX1 \recentABools_len_reg[7]  ( .D(n4333), .CLK(n9139), .Q(
        recentABools_len[7]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[8]  ( .D(n4268), .CLK(n9139), .Q(
        recentABools_len_new_reg_385[8]) );
  DFFPOSX1 \recentABools_len_reg[8]  ( .D(n4332), .CLK(n9139), .Q(
        recentABools_len[8]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[9]  ( .D(n4267), .CLK(n9139), .Q(
        recentABools_len_new_reg_385[9]) );
  DFFPOSX1 \recentABools_len_reg[9]  ( .D(n4331), .CLK(n9139), .Q(
        recentABools_len[9]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[10]  ( .D(n4266), .CLK(n9139), 
        .Q(recentABools_len_new_reg_385[10]) );
  DFFPOSX1 \recentABools_len_reg[10]  ( .D(n4330), .CLK(n9139), .Q(
        recentABools_len[10]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[11]  ( .D(n4265), .CLK(n9138), 
        .Q(recentABools_len_new_reg_385[11]) );
  DFFPOSX1 \recentABools_len_reg[11]  ( .D(n4329), .CLK(n9138), .Q(
        recentABools_len[11]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[12]  ( .D(n4264), .CLK(n9138), 
        .Q(recentABools_len_new_reg_385[12]) );
  DFFPOSX1 \recentABools_len_reg[12]  ( .D(n4328), .CLK(n9138), .Q(
        recentABools_len[12]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[13]  ( .D(n4263), .CLK(n9138), 
        .Q(recentABools_len_new_reg_385[13]) );
  DFFPOSX1 \recentABools_len_reg[13]  ( .D(n4327), .CLK(n9138), .Q(
        recentABools_len[13]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[14]  ( .D(n4262), .CLK(n9138), 
        .Q(recentABools_len_new_reg_385[14]) );
  DFFPOSX1 \recentABools_len_reg[14]  ( .D(n4326), .CLK(n9138), .Q(
        recentABools_len[14]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[15]  ( .D(n4261), .CLK(n9138), 
        .Q(recentABools_len_new_reg_385[15]) );
  DFFPOSX1 \recentABools_len_reg[15]  ( .D(n4325), .CLK(n9138), .Q(
        recentABools_len[15]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[16]  ( .D(n4260), .CLK(n9138), 
        .Q(recentABools_len_new_reg_385[16]) );
  DFFPOSX1 \recentABools_len_reg[16]  ( .D(n4324), .CLK(n9138), .Q(
        recentABools_len[16]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[17]  ( .D(n4259), .CLK(n9138), 
        .Q(recentABools_len_new_reg_385[17]) );
  DFFPOSX1 \recentABools_len_reg[17]  ( .D(n4323), .CLK(n9137), .Q(
        recentABools_len[17]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[18]  ( .D(n4258), .CLK(n9137), 
        .Q(recentABools_len_new_reg_385[18]) );
  DFFPOSX1 \recentABools_len_reg[18]  ( .D(n4322), .CLK(n9137), .Q(
        recentABools_len[18]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[19]  ( .D(n4257), .CLK(n9137), 
        .Q(recentABools_len_new_reg_385[19]) );
  DFFPOSX1 \recentABools_len_reg[19]  ( .D(n4321), .CLK(n9137), .Q(
        recentABools_len[19]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[20]  ( .D(n4256), .CLK(n9137), 
        .Q(recentABools_len_new_reg_385[20]) );
  DFFPOSX1 \recentABools_len_reg[20]  ( .D(n4320), .CLK(n9137), .Q(
        recentABools_len[20]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[21]  ( .D(n4255), .CLK(n9137), 
        .Q(recentABools_len_new_reg_385[21]) );
  DFFPOSX1 \recentABools_len_reg[21]  ( .D(n4319), .CLK(n9137), .Q(
        recentABools_len[21]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[22]  ( .D(n4254), .CLK(n9137), 
        .Q(recentABools_len_new_reg_385[22]) );
  DFFPOSX1 \recentABools_len_reg[22]  ( .D(n4318), .CLK(n9137), .Q(
        recentABools_len[22]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[23]  ( .D(n4253), .CLK(n9137), 
        .Q(recentABools_len_new_reg_385[23]) );
  DFFPOSX1 \recentABools_len_reg[23]  ( .D(n4317), .CLK(n9137), .Q(
        recentABools_len[23]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[24]  ( .D(n4252), .CLK(n9136), 
        .Q(recentABools_len_new_reg_385[24]) );
  DFFPOSX1 \recentABools_len_reg[24]  ( .D(n4316), .CLK(n9136), .Q(
        recentABools_len[24]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[25]  ( .D(n4251), .CLK(n9136), 
        .Q(recentABools_len_new_reg_385[25]) );
  DFFPOSX1 \recentABools_len_reg[25]  ( .D(n4315), .CLK(n9136), .Q(
        recentABools_len[25]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[26]  ( .D(n4250), .CLK(n9136), 
        .Q(recentABools_len_new_reg_385[26]) );
  DFFPOSX1 \recentABools_len_reg[26]  ( .D(n4314), .CLK(n9136), .Q(
        recentABools_len[26]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[27]  ( .D(n4249), .CLK(n9136), 
        .Q(recentABools_len_new_reg_385[27]) );
  DFFPOSX1 \recentABools_len_reg[27]  ( .D(n4313), .CLK(n9136), .Q(
        recentABools_len[27]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[28]  ( .D(n4248), .CLK(n9136), 
        .Q(recentABools_len_new_reg_385[28]) );
  DFFPOSX1 \recentABools_len_reg[28]  ( .D(n4312), .CLK(n9136), .Q(
        recentABools_len[28]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[29]  ( .D(n4247), .CLK(n9136), 
        .Q(recentABools_len_new_reg_385[29]) );
  DFFPOSX1 \recentABools_len_reg[29]  ( .D(n4311), .CLK(n9136), .Q(
        recentABools_len[29]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[0]  ( .D(n3486), 
        .CLK(n9136), .Q(CircularBuffer_len_write_assig_2_reg_1729[0]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[1]  ( .D(n3485), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[1]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[2]  ( .D(n3484), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[2]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[3]  ( .D(n3483), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[3]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[4]  ( .D(n3482), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[4]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[5]  ( .D(n3481), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[5]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[6]  ( .D(n3480), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[6]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[7]  ( .D(n3479), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[7]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[8]  ( .D(n3478), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[8]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[9]  ( .D(n3477), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[9]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[10]  ( .D(n3476), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[10]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[11]  ( .D(n3475), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[11]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[12]  ( .D(n3474), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[12]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[13]  ( .D(n3473), 
        .CLK(n9135), .Q(CircularBuffer_len_write_assig_2_reg_1729[13]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[14]  ( .D(n3472), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[14]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[15]  ( .D(n3471), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[15]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[16]  ( .D(n3470), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[16]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[17]  ( .D(n3469), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[17]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[18]  ( .D(n3468), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[18]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[19]  ( .D(n3467), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[19]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[20]  ( .D(n3466), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[20]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[21]  ( .D(n3465), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[21]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[22]  ( .D(n3464), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[22]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[23]  ( .D(n3463), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[23]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[24]  ( .D(n3462), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[24]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[25]  ( .D(n3461), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[25]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[26]  ( .D(n3460), 
        .CLK(n9134), .Q(CircularBuffer_len_write_assig_2_reg_1729[26]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[27]  ( .D(n3459), 
        .CLK(n9133), .Q(CircularBuffer_len_write_assig_2_reg_1729[27]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[28]  ( .D(n3458), 
        .CLK(n9133), .Q(CircularBuffer_len_write_assig_2_reg_1729[28]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[29]  ( .D(n3457), 
        .CLK(n9133), .Q(CircularBuffer_len_write_assig_2_reg_1729[29]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[30]  ( .D(n3456), 
        .CLK(n9133), .Q(CircularBuffer_len_write_assig_2_reg_1729[30]) );
  DFFPOSX1 \CircularBuffer_len_write_assig_2_reg_1729_reg[31]  ( .D(n3455), 
        .CLK(n9133), .Q(CircularBuffer_len_write_assig_2_reg_1729[31]) );
  DFFPOSX1 \recentABools_data_load_reg_1700_reg[0]  ( .D(n3454), .CLK(n9133), 
        .Q(\recentABools_data_load_reg_1700[0] ) );
  DFFPOSX1 \toReturn_7_reg_1750_reg[0]  ( .D(n3453), .CLK(n9133), .Q(
        \toReturn_7_reg_1750[0] ) );
  DFFPOSX1 \not_tmp_i_i2_reg_1745_reg[0]  ( .D(n4717), .CLK(n9133), .Q(
        \not_tmp_i_i2_reg_1745[0] ) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[31]  ( .D(n4341), .CLK(n9133), 
        .Q(recentABools_len_new_reg_385[31]) );
  DFFPOSX1 \recentABools_len_reg[31]  ( .D(n4309), .CLK(n9133), .Q(
        recentABools_len[31]) );
  DFFPOSX1 \recentABools_len_new_reg_385_reg[0]  ( .D(n4276), .CLK(n9133), .Q(
        recentABools_len_new_reg_385[0]) );
  DFFPOSX1 \ap_CS_fsm_reg[13]  ( .D(N111), .CLK(n9133), .Q(ap_CS_fsm[13]) );
  DFFPOSX1 \AbeatDelay_reg[0]  ( .D(n3451), .CLK(n9133), .Q(AbeatDelay[0]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[0]  ( .D(n3450), .CLK(n9132), .Q(
        tmp_3_reg_1589[0]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[0]  ( .D(n4244), .CLK(n9132), .Q(
        AbeatDelay_new_reg_394[0]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[1]  ( .D(n3449), .CLK(n9132), .Q(
        tmp_3_reg_1589[1]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[1]  ( .D(n4243), .CLK(n9132), .Q(
        AbeatDelay_new_reg_394[1]) );
  DFFPOSX1 \AbeatDelay_reg[1]  ( .D(n3448), .CLK(n9132), .Q(AbeatDelay[1]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[2]  ( .D(n3447), .CLK(n9132), .Q(
        tmp_3_reg_1589[2]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[2]  ( .D(n4242), .CLK(n9132), .Q(
        AbeatDelay_new_reg_394[2]) );
  DFFPOSX1 \AbeatDelay_reg[2]  ( .D(n3446), .CLK(n9132), .Q(AbeatDelay[2]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[3]  ( .D(n3445), .CLK(n9132), .Q(
        tmp_3_reg_1589[3]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[3]  ( .D(n4241), .CLK(n9132), .Q(
        AbeatDelay_new_reg_394[3]) );
  DFFPOSX1 \AbeatDelay_reg[3]  ( .D(n3444), .CLK(n9132), .Q(AbeatDelay[3]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[4]  ( .D(n3443), .CLK(n9132), .Q(
        tmp_3_reg_1589[4]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[4]  ( .D(n4240), .CLK(n9132), .Q(
        AbeatDelay_new_reg_394[4]) );
  DFFPOSX1 \AbeatDelay_reg[4]  ( .D(n3442), .CLK(n9131), .Q(AbeatDelay[4]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[5]  ( .D(n3441), .CLK(n9131), .Q(
        tmp_3_reg_1589[5]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[5]  ( .D(n4239), .CLK(n9131), .Q(
        AbeatDelay_new_reg_394[5]) );
  DFFPOSX1 \AbeatDelay_reg[5]  ( .D(n3440), .CLK(n9131), .Q(AbeatDelay[5]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[6]  ( .D(n3439), .CLK(n9131), .Q(
        tmp_3_reg_1589[6]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[6]  ( .D(n4238), .CLK(n9131), .Q(
        AbeatDelay_new_reg_394[6]) );
  DFFPOSX1 \AbeatDelay_reg[6]  ( .D(n3438), .CLK(n9131), .Q(AbeatDelay[6]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[7]  ( .D(n3437), .CLK(n9131), .Q(
        tmp_3_reg_1589[7]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[7]  ( .D(n4237), .CLK(n9131), .Q(
        AbeatDelay_new_reg_394[7]) );
  DFFPOSX1 \AbeatDelay_reg[7]  ( .D(n3436), .CLK(n9131), .Q(AbeatDelay[7]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[8]  ( .D(n3435), .CLK(n9131), .Q(
        tmp_3_reg_1589[8]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[8]  ( .D(n4236), .CLK(n9131), .Q(
        AbeatDelay_new_reg_394[8]) );
  DFFPOSX1 \AbeatDelay_reg[8]  ( .D(n3434), .CLK(n9131), .Q(AbeatDelay[8]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[9]  ( .D(n3433), .CLK(n9130), .Q(
        tmp_3_reg_1589[9]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[9]  ( .D(n4235), .CLK(n9130), .Q(
        AbeatDelay_new_reg_394[9]) );
  DFFPOSX1 \AbeatDelay_reg[9]  ( .D(n3432), .CLK(n9130), .Q(AbeatDelay[9]) );
  DFFPOSX1 \tmp_3_reg_1589_reg[10]  ( .D(n3431), .CLK(n9130), .Q(
        tmp_3_reg_1589[10]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[10]  ( .D(n4234), .CLK(n9130), .Q(
        AbeatDelay_new_reg_394[10]) );
  DFFPOSX1 \AbeatDelay_reg[10]  ( .D(n3430), .CLK(n9130), .Q(AbeatDelay[10])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[11]  ( .D(n3429), .CLK(n9130), .Q(
        tmp_3_reg_1589[11]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[11]  ( .D(n4233), .CLK(n9130), .Q(
        AbeatDelay_new_reg_394[11]) );
  DFFPOSX1 \AbeatDelay_reg[11]  ( .D(n3428), .CLK(n9130), .Q(AbeatDelay[11])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[12]  ( .D(n3427), .CLK(n9130), .Q(
        tmp_3_reg_1589[12]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[12]  ( .D(n4232), .CLK(n9130), .Q(
        AbeatDelay_new_reg_394[12]) );
  DFFPOSX1 \AbeatDelay_reg[12]  ( .D(n3426), .CLK(n9130), .Q(AbeatDelay[12])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[13]  ( .D(n3425), .CLK(n9130), .Q(
        tmp_3_reg_1589[13]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[13]  ( .D(n4231), .CLK(n9129), .Q(
        AbeatDelay_new_reg_394[13]) );
  DFFPOSX1 \AbeatDelay_reg[13]  ( .D(n3424), .CLK(n9129), .Q(AbeatDelay[13])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[14]  ( .D(n3423), .CLK(n9129), .Q(
        tmp_3_reg_1589[14]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[14]  ( .D(n4230), .CLK(n9129), .Q(
        AbeatDelay_new_reg_394[14]) );
  DFFPOSX1 \AbeatDelay_reg[14]  ( .D(n3422), .CLK(n9129), .Q(AbeatDelay[14])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[15]  ( .D(n3421), .CLK(n9129), .Q(
        tmp_3_reg_1589[15]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[15]  ( .D(n4229), .CLK(n9129), .Q(
        AbeatDelay_new_reg_394[15]) );
  DFFPOSX1 \AbeatDelay_reg[15]  ( .D(n3420), .CLK(n9129), .Q(AbeatDelay[15])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[16]  ( .D(n3419), .CLK(n9129), .Q(
        tmp_3_reg_1589[16]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[16]  ( .D(n4228), .CLK(n9129), .Q(
        AbeatDelay_new_reg_394[16]) );
  DFFPOSX1 \AbeatDelay_reg[16]  ( .D(n3418), .CLK(n9129), .Q(AbeatDelay[16])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[17]  ( .D(n3417), .CLK(n9129), .Q(
        tmp_3_reg_1589[17]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[17]  ( .D(n4227), .CLK(n9129), .Q(
        AbeatDelay_new_reg_394[17]) );
  DFFPOSX1 \AbeatDelay_reg[17]  ( .D(n3416), .CLK(n9128), .Q(AbeatDelay[17])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[18]  ( .D(n3415), .CLK(n9128), .Q(
        tmp_3_reg_1589[18]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[18]  ( .D(n4226), .CLK(n9128), .Q(
        AbeatDelay_new_reg_394[18]) );
  DFFPOSX1 \AbeatDelay_reg[18]  ( .D(n3414), .CLK(n9128), .Q(AbeatDelay[18])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[19]  ( .D(n3413), .CLK(n9128), .Q(
        tmp_3_reg_1589[19]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[19]  ( .D(n4225), .CLK(n9128), .Q(
        AbeatDelay_new_reg_394[19]) );
  DFFPOSX1 \AbeatDelay_reg[19]  ( .D(n3412), .CLK(n9128), .Q(AbeatDelay[19])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[20]  ( .D(n3411), .CLK(n9128), .Q(
        tmp_3_reg_1589[20]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[20]  ( .D(n4224), .CLK(n9128), .Q(
        AbeatDelay_new_reg_394[20]) );
  DFFPOSX1 \AbeatDelay_reg[20]  ( .D(n3410), .CLK(n9128), .Q(AbeatDelay[20])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[21]  ( .D(n3409), .CLK(n9128), .Q(
        tmp_3_reg_1589[21]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[21]  ( .D(n4223), .CLK(n9128), .Q(
        AbeatDelay_new_reg_394[21]) );
  DFFPOSX1 \AbeatDelay_reg[21]  ( .D(n3408), .CLK(n9128), .Q(AbeatDelay[21])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[22]  ( .D(n3407), .CLK(n9127), .Q(
        tmp_3_reg_1589[22]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[22]  ( .D(n4222), .CLK(n9127), .Q(
        AbeatDelay_new_reg_394[22]) );
  DFFPOSX1 \AbeatDelay_reg[22]  ( .D(n3406), .CLK(n9127), .Q(AbeatDelay[22])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[23]  ( .D(n3405), .CLK(n9127), .Q(
        tmp_3_reg_1589[23]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[23]  ( .D(n4221), .CLK(n9127), .Q(
        AbeatDelay_new_reg_394[23]) );
  DFFPOSX1 \AbeatDelay_reg[23]  ( .D(n3404), .CLK(n9127), .Q(AbeatDelay[23])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[24]  ( .D(n3403), .CLK(n9127), .Q(
        tmp_3_reg_1589[24]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[24]  ( .D(n4220), .CLK(n9127), .Q(
        AbeatDelay_new_reg_394[24]) );
  DFFPOSX1 \AbeatDelay_reg[24]  ( .D(n3402), .CLK(n9127), .Q(AbeatDelay[24])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[25]  ( .D(n3401), .CLK(n9127), .Q(
        tmp_3_reg_1589[25]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[25]  ( .D(n4219), .CLK(n9127), .Q(
        AbeatDelay_new_reg_394[25]) );
  DFFPOSX1 \AbeatDelay_reg[25]  ( .D(n3400), .CLK(n9127), .Q(AbeatDelay[25])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[26]  ( .D(n3399), .CLK(n9127), .Q(
        tmp_3_reg_1589[26]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[26]  ( .D(n4218), .CLK(n9126), .Q(
        AbeatDelay_new_reg_394[26]) );
  DFFPOSX1 \AbeatDelay_reg[26]  ( .D(n3398), .CLK(n9126), .Q(AbeatDelay[26])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[27]  ( .D(n3397), .CLK(n9126), .Q(
        tmp_3_reg_1589[27]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[27]  ( .D(n4217), .CLK(n9126), .Q(
        AbeatDelay_new_reg_394[27]) );
  DFFPOSX1 \AbeatDelay_reg[27]  ( .D(n3396), .CLK(n9126), .Q(AbeatDelay[27])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[28]  ( .D(n3395), .CLK(n9126), .Q(
        tmp_3_reg_1589[28]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[28]  ( .D(n4216), .CLK(n9126), .Q(
        AbeatDelay_new_reg_394[28]) );
  DFFPOSX1 \AbeatDelay_reg[28]  ( .D(n3394), .CLK(n9126), .Q(AbeatDelay[28])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[29]  ( .D(n3393), .CLK(n9126), .Q(
        tmp_3_reg_1589[29]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[29]  ( .D(n4215), .CLK(n9126), .Q(
        AbeatDelay_new_reg_394[29]) );
  DFFPOSX1 \AbeatDelay_reg[29]  ( .D(n3392), .CLK(n9126), .Q(AbeatDelay[29])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[30]  ( .D(n3391), .CLK(n9126), .Q(
        tmp_3_reg_1589[30]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[30]  ( .D(n4214), .CLK(n9126), .Q(
        AbeatDelay_new_reg_394[30]) );
  DFFPOSX1 \AbeatDelay_reg[30]  ( .D(n3390), .CLK(n9125), .Q(AbeatDelay[30])
         );
  DFFPOSX1 \tmp_3_reg_1589_reg[31]  ( .D(n3389), .CLK(n9125), .Q(
        tmp_3_reg_1589[31]) );
  DFFPOSX1 \AbeatDelay_new_reg_394_reg[31]  ( .D(n4680), .CLK(n9125), .Q(
        AbeatDelay_new_reg_394[31]) );
  DFFPOSX1 \AbeatDelay_reg[31]  ( .D(n3388), .CLK(n9125), .Q(AbeatDelay[31])
         );
  DFFPOSX1 \AstimDelay_reg[0]  ( .D(n3387), .CLK(n9125), .Q(AstimDelay[0]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[0]  ( .D(n3386), .CLK(n9125), .Q(
        tmp_6_reg_1538[0]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[1]  ( .D(n3385), .CLK(n9125), .Q(
        tmp_6_reg_1538[1]) );
  DFFPOSX1 \AstimDelay_reg[1]  ( .D(n3384), .CLK(n9125), .Q(AstimDelay[1]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[2]  ( .D(n3383), .CLK(n9125), .Q(
        tmp_6_reg_1538[2]) );
  DFFPOSX1 \AstimDelay_reg[2]  ( .D(n3382), .CLK(n9125), .Q(AstimDelay[2]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[3]  ( .D(n3381), .CLK(n9125), .Q(
        tmp_6_reg_1538[3]) );
  DFFPOSX1 \AstimDelay_reg[3]  ( .D(n3380), .CLK(n9125), .Q(AstimDelay[3]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[4]  ( .D(n3379), .CLK(n9125), .Q(
        tmp_6_reg_1538[4]) );
  DFFPOSX1 \AstimDelay_reg[4]  ( .D(n3378), .CLK(n9124), .Q(AstimDelay[4]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[5]  ( .D(n3377), .CLK(n9124), .Q(
        tmp_6_reg_1538[5]) );
  DFFPOSX1 \AstimDelay_reg[5]  ( .D(n3376), .CLK(n9124), .Q(AstimDelay[5]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[6]  ( .D(n3375), .CLK(n9124), .Q(
        tmp_6_reg_1538[6]) );
  DFFPOSX1 \AstimDelay_reg[6]  ( .D(n3374), .CLK(n9124), .Q(AstimDelay[6]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[7]  ( .D(n3373), .CLK(n9124), .Q(
        tmp_6_reg_1538[7]) );
  DFFPOSX1 \AstimDelay_reg[7]  ( .D(n3372), .CLK(n9124), .Q(AstimDelay[7]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[8]  ( .D(n3371), .CLK(n9124), .Q(
        tmp_6_reg_1538[8]) );
  DFFPOSX1 \AstimDelay_reg[8]  ( .D(n3370), .CLK(n9124), .Q(AstimDelay[8]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[9]  ( .D(n3369), .CLK(n9124), .Q(
        tmp_6_reg_1538[9]) );
  DFFPOSX1 \AstimDelay_reg[9]  ( .D(n3368), .CLK(n9124), .Q(AstimDelay[9]) );
  DFFPOSX1 \tmp_6_reg_1538_reg[10]  ( .D(n3367), .CLK(n9124), .Q(
        tmp_6_reg_1538[10]) );
  DFFPOSX1 \AstimDelay_reg[10]  ( .D(n3366), .CLK(n9124), .Q(AstimDelay[10])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[11]  ( .D(n3365), .CLK(n9123), .Q(
        tmp_6_reg_1538[11]) );
  DFFPOSX1 \AstimDelay_reg[11]  ( .D(n3364), .CLK(n9123), .Q(AstimDelay[11])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[12]  ( .D(n3363), .CLK(n9123), .Q(
        tmp_6_reg_1538[12]) );
  DFFPOSX1 \AstimDelay_reg[12]  ( .D(n3362), .CLK(n9123), .Q(AstimDelay[12])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[13]  ( .D(n3361), .CLK(n9123), .Q(
        tmp_6_reg_1538[13]) );
  DFFPOSX1 \AstimDelay_reg[13]  ( .D(n3360), .CLK(n9123), .Q(AstimDelay[13])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[14]  ( .D(n3359), .CLK(n9123), .Q(
        tmp_6_reg_1538[14]) );
  DFFPOSX1 \AstimDelay_reg[14]  ( .D(n3358), .CLK(n9123), .Q(AstimDelay[14])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[15]  ( .D(n3357), .CLK(n9123), .Q(
        tmp_6_reg_1538[15]) );
  DFFPOSX1 \AstimDelay_reg[15]  ( .D(n3356), .CLK(n9123), .Q(AstimDelay[15])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[16]  ( .D(n3355), .CLK(n9123), .Q(
        tmp_6_reg_1538[16]) );
  DFFPOSX1 \AstimDelay_reg[16]  ( .D(n3354), .CLK(n9123), .Q(AstimDelay[16])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[17]  ( .D(n3353), .CLK(n9123), .Q(
        tmp_6_reg_1538[17]) );
  DFFPOSX1 \AstimDelay_reg[17]  ( .D(n3352), .CLK(n9122), .Q(AstimDelay[17])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[18]  ( .D(n3351), .CLK(n9122), .Q(
        tmp_6_reg_1538[18]) );
  DFFPOSX1 \AstimDelay_reg[18]  ( .D(n3350), .CLK(n9122), .Q(AstimDelay[18])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[19]  ( .D(n3349), .CLK(n9122), .Q(
        tmp_6_reg_1538[19]) );
  DFFPOSX1 \AstimDelay_reg[19]  ( .D(n3348), .CLK(n9122), .Q(AstimDelay[19])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[20]  ( .D(n3347), .CLK(n9122), .Q(
        tmp_6_reg_1538[20]) );
  DFFPOSX1 \AstimDelay_reg[20]  ( .D(n3346), .CLK(n9122), .Q(AstimDelay[20])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[21]  ( .D(n3345), .CLK(n9122), .Q(
        tmp_6_reg_1538[21]) );
  DFFPOSX1 \AstimDelay_reg[21]  ( .D(n3344), .CLK(n9122), .Q(AstimDelay[21])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[22]  ( .D(n3343), .CLK(n9122), .Q(
        tmp_6_reg_1538[22]) );
  DFFPOSX1 \AstimDelay_reg[22]  ( .D(n3342), .CLK(n9122), .Q(AstimDelay[22])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[23]  ( .D(n3341), .CLK(n9122), .Q(
        tmp_6_reg_1538[23]) );
  DFFPOSX1 \AstimDelay_reg[23]  ( .D(n3340), .CLK(n9122), .Q(AstimDelay[23])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[24]  ( .D(n3339), .CLK(n9121), .Q(
        tmp_6_reg_1538[24]) );
  DFFPOSX1 \AstimDelay_reg[24]  ( .D(n3338), .CLK(n9121), .Q(AstimDelay[24])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[25]  ( .D(n3337), .CLK(n9121), .Q(
        tmp_6_reg_1538[25]) );
  DFFPOSX1 \AstimDelay_reg[25]  ( .D(n3336), .CLK(n9121), .Q(AstimDelay[25])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[26]  ( .D(n3335), .CLK(n9121), .Q(
        tmp_6_reg_1538[26]) );
  DFFPOSX1 \AstimDelay_reg[26]  ( .D(n3334), .CLK(n9121), .Q(AstimDelay[26])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[27]  ( .D(n3333), .CLK(n9121), .Q(
        tmp_6_reg_1538[27]) );
  DFFPOSX1 \AstimDelay_reg[27]  ( .D(n3332), .CLK(n9121), .Q(AstimDelay[27])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[28]  ( .D(n3331), .CLK(n9121), .Q(
        tmp_6_reg_1538[28]) );
  DFFPOSX1 \AstimDelay_reg[28]  ( .D(n3330), .CLK(n9121), .Q(AstimDelay[28])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[29]  ( .D(n3329), .CLK(n9121), .Q(
        tmp_6_reg_1538[29]) );
  DFFPOSX1 \AstimDelay_reg[29]  ( .D(n3328), .CLK(n9121), .Q(AstimDelay[29])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[30]  ( .D(n3327), .CLK(n9121), .Q(
        tmp_6_reg_1538[30]) );
  DFFPOSX1 \AstimDelay_reg[30]  ( .D(n3326), .CLK(n9120), .Q(AstimDelay[30])
         );
  DFFPOSX1 \tmp_6_reg_1538_reg[31]  ( .D(n3325), .CLK(n9120), .Q(
        tmp_6_reg_1538[31]) );
  DFFPOSX1 \tmp_22_reg_1772_reg[0]  ( .D(n3324), .CLK(n9120), .Q(
        \tmp_22_reg_1772[0] ) );
  DFFPOSX1 \AstimDelay_reg[31]  ( .D(n3323), .CLK(n9120), .Q(AstimDelay[31])
         );
  DFFPOSX1 \VstimDelay_reg[0]  ( .D(n3322), .CLK(n9120), .Q(VstimDelay[0]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[0]  ( .D(n3321), .CLK(n9120), .Q(
        tmp_7_reg_1544[0]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[1]  ( .D(n3320), .CLK(n9120), .Q(
        tmp_7_reg_1544[1]) );
  DFFPOSX1 \VstimDelay_reg[1]  ( .D(n3319), .CLK(n9120), .Q(VstimDelay[1]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[2]  ( .D(n3318), .CLK(n9120), .Q(
        tmp_7_reg_1544[2]) );
  DFFPOSX1 \VstimDelay_reg[2]  ( .D(n3317), .CLK(n9120), .Q(VstimDelay[2]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[3]  ( .D(n3316), .CLK(n9120), .Q(
        tmp_7_reg_1544[3]) );
  DFFPOSX1 \VstimDelay_reg[3]  ( .D(n3315), .CLK(n9120), .Q(VstimDelay[3]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[4]  ( .D(n3314), .CLK(n9120), .Q(
        tmp_7_reg_1544[4]) );
  DFFPOSX1 \VstimDelay_reg[4]  ( .D(n3313), .CLK(n9119), .Q(VstimDelay[4]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[5]  ( .D(n3312), .CLK(n9119), .Q(
        tmp_7_reg_1544[5]) );
  DFFPOSX1 \VstimDelay_reg[5]  ( .D(n3311), .CLK(n9119), .Q(VstimDelay[5]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[6]  ( .D(n3310), .CLK(n9119), .Q(
        tmp_7_reg_1544[6]) );
  DFFPOSX1 \VstimDelay_reg[6]  ( .D(n3309), .CLK(n9119), .Q(VstimDelay[6]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[7]  ( .D(n3308), .CLK(n9119), .Q(
        tmp_7_reg_1544[7]) );
  DFFPOSX1 \VstimDelay_reg[7]  ( .D(n3307), .CLK(n9119), .Q(VstimDelay[7]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[8]  ( .D(n3306), .CLK(n9119), .Q(
        tmp_7_reg_1544[8]) );
  DFFPOSX1 \VstimDelay_reg[8]  ( .D(n3305), .CLK(n9119), .Q(VstimDelay[8]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[9]  ( .D(n3304), .CLK(n9119), .Q(
        tmp_7_reg_1544[9]) );
  DFFPOSX1 \VstimDelay_reg[9]  ( .D(n3303), .CLK(n9119), .Q(VstimDelay[9]) );
  DFFPOSX1 \tmp_7_reg_1544_reg[10]  ( .D(n3302), .CLK(n9119), .Q(
        tmp_7_reg_1544[10]) );
  DFFPOSX1 \VstimDelay_reg[10]  ( .D(n3301), .CLK(n9119), .Q(VstimDelay[10])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[11]  ( .D(n3300), .CLK(n9118), .Q(
        tmp_7_reg_1544[11]) );
  DFFPOSX1 \VstimDelay_reg[11]  ( .D(n3299), .CLK(n9118), .Q(VstimDelay[11])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[12]  ( .D(n3298), .CLK(n9118), .Q(
        tmp_7_reg_1544[12]) );
  DFFPOSX1 \VstimDelay_reg[12]  ( .D(n3297), .CLK(n9118), .Q(VstimDelay[12])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[13]  ( .D(n3296), .CLK(n9118), .Q(
        tmp_7_reg_1544[13]) );
  DFFPOSX1 \VstimDelay_reg[13]  ( .D(n3295), .CLK(n9118), .Q(VstimDelay[13])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[14]  ( .D(n3294), .CLK(n9118), .Q(
        tmp_7_reg_1544[14]) );
  DFFPOSX1 \VstimDelay_reg[14]  ( .D(n3293), .CLK(n9118), .Q(VstimDelay[14])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[15]  ( .D(n3292), .CLK(n9118), .Q(
        tmp_7_reg_1544[15]) );
  DFFPOSX1 \VstimDelay_reg[15]  ( .D(n3291), .CLK(n9118), .Q(VstimDelay[15])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[16]  ( .D(n3290), .CLK(n9118), .Q(
        tmp_7_reg_1544[16]) );
  DFFPOSX1 \VstimDelay_reg[16]  ( .D(n3289), .CLK(n9118), .Q(VstimDelay[16])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[17]  ( .D(n3288), .CLK(n9118), .Q(
        tmp_7_reg_1544[17]) );
  DFFPOSX1 \VstimDelay_reg[17]  ( .D(n3287), .CLK(n9117), .Q(VstimDelay[17])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[18]  ( .D(n3286), .CLK(n9117), .Q(
        tmp_7_reg_1544[18]) );
  DFFPOSX1 \VstimDelay_reg[18]  ( .D(n3285), .CLK(n9117), .Q(VstimDelay[18])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[19]  ( .D(n3284), .CLK(n9117), .Q(
        tmp_7_reg_1544[19]) );
  DFFPOSX1 \VstimDelay_reg[19]  ( .D(n3283), .CLK(n9117), .Q(VstimDelay[19])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[20]  ( .D(n3282), .CLK(n9117), .Q(
        tmp_7_reg_1544[20]) );
  DFFPOSX1 \VstimDelay_reg[20]  ( .D(n3281), .CLK(n9117), .Q(VstimDelay[20])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[21]  ( .D(n3280), .CLK(n9117), .Q(
        tmp_7_reg_1544[21]) );
  DFFPOSX1 \VstimDelay_reg[21]  ( .D(n3279), .CLK(n9117), .Q(VstimDelay[21])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[22]  ( .D(n3278), .CLK(n9117), .Q(
        tmp_7_reg_1544[22]) );
  DFFPOSX1 \VstimDelay_reg[22]  ( .D(n3277), .CLK(n9117), .Q(VstimDelay[22])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[23]  ( .D(n3276), .CLK(n9117), .Q(
        tmp_7_reg_1544[23]) );
  DFFPOSX1 \VstimDelay_reg[23]  ( .D(n3275), .CLK(n9117), .Q(VstimDelay[23])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[24]  ( .D(n3274), .CLK(n9116), .Q(
        tmp_7_reg_1544[24]) );
  DFFPOSX1 \VstimDelay_reg[24]  ( .D(n3273), .CLK(n9116), .Q(VstimDelay[24])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[25]  ( .D(n3272), .CLK(n9116), .Q(
        tmp_7_reg_1544[25]) );
  DFFPOSX1 \VstimDelay_reg[25]  ( .D(n3271), .CLK(n9116), .Q(VstimDelay[25])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[26]  ( .D(n3270), .CLK(n9116), .Q(
        tmp_7_reg_1544[26]) );
  DFFPOSX1 \VstimDelay_reg[26]  ( .D(n3269), .CLK(n9116), .Q(VstimDelay[26])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[27]  ( .D(n3268), .CLK(n9116), .Q(
        tmp_7_reg_1544[27]) );
  DFFPOSX1 \VstimDelay_reg[27]  ( .D(n3267), .CLK(n9116), .Q(VstimDelay[27])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[28]  ( .D(n3266), .CLK(n9116), .Q(
        tmp_7_reg_1544[28]) );
  DFFPOSX1 \VstimDelay_reg[28]  ( .D(n3265), .CLK(n9116), .Q(VstimDelay[28])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[29]  ( .D(n3264), .CLK(n9116), .Q(
        tmp_7_reg_1544[29]) );
  DFFPOSX1 \VstimDelay_reg[29]  ( .D(n3263), .CLK(n9116), .Q(VstimDelay[29])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[30]  ( .D(n3262), .CLK(n9116), .Q(
        tmp_7_reg_1544[30]) );
  DFFPOSX1 \VstimDelay_reg[30]  ( .D(n3261), .CLK(n9115), .Q(VstimDelay[30])
         );
  DFFPOSX1 \tmp_7_reg_1544_reg[31]  ( .D(n3260), .CLK(n9115), .Q(
        tmp_7_reg_1544[31]) );
  DFFPOSX1 \tmp_25_reg_1777_reg[0]  ( .D(n3259), .CLK(n9115), .Q(
        \tmp_25_reg_1777[0] ) );
  DFFPOSX1 \VstimDelay_reg[31]  ( .D(n3258), .CLK(n9115), .Q(VstimDelay[31])
         );
  DFFPOSX1 \last_sample_is_A_V_reg[0]  ( .D(n4245), .CLK(n9115), .Q(
        \last_sample_is_A_V[0] ) );
  DFFPOSX1 \recentABools_sum_reg[30]  ( .D(n4372), .CLK(n9115), .Q(
        recentABools_sum[30]) );
  DFFPOSX1 \CircularBuffer_sum_read_assign_1_reg_1705_reg[31]  ( .D(n3257), 
        .CLK(n9115), .Q(CircularBuffer_sum_read_assign_1_reg_1705[31]) );
  DFFPOSX1 \sum_1_reg_376_reg[31]  ( .D(n4277), .CLK(n9115), .Q(
        sum_1_reg_376[31]) );
  NOR3X1 U3 ( .A(n5897), .B(n5901), .C(n5907), .Y(toReturn_1_fu_1395_p3_12) );
  NOR3X1 U5 ( .A(n7602), .B(AbeatDelay_new_reg_394[12]), .C(
        AbeatDelay_new_reg_394[11]), .Y(n268) );
  NOR3X1 U7 ( .A(n7415), .B(n8393), .C(n9385), .Y(n267) );
  NOR3X1 U10 ( .A(n7085), .B(AbeatDelay_new_reg_394[1]), .C(
        AbeatDelay_new_reg_394[19]), .Y(n277) );
  NAND3X1 U11 ( .A(n10721), .B(n10723), .C(n10719), .Y(n278) );
  NOR3X1 U12 ( .A(n7244), .B(AbeatDelay_new_reg_394[16]), .C(
        AbeatDelay_new_reg_394[15]), .Y(n276) );
  NAND3X1 U14 ( .A(n285), .B(n286), .C(n287), .Y(n264) );
  NOR3X1 U15 ( .A(n5896), .B(n5900), .C(n5906), .Y(n287) );
  NAND3X1 U17 ( .A(n10695), .B(n10697), .C(n10693), .Y(n289) );
  NAND3X1 U18 ( .A(n10739), .B(n10741), .C(n8265), .Y(n288) );
  NOR3X1 U20 ( .A(n8282), .B(AbeatDelay_new_reg_394[28]), .C(
        AbeatDelay_new_reg_394[27]), .Y(n286) );
  NOR3X1 U22 ( .A(n7801), .B(AbeatDelay_new_reg_394[24]), .C(
        AbeatDelay_new_reg_394[23]), .Y(n285) );
  NAND3X1 U25 ( .A(n307), .B(n308), .C(n309), .Y(n306) );
  NOR3X1 U26 ( .A(n7815), .B(n7813), .C(n7814), .Y(n309) );
  NAND3X1 U33 ( .A(\last_sample_is_V_V_loc_2_reg_358[0] ), .B(n10451), .C(
        n8014), .Y(n310) );
  NOR3X1 U35 ( .A(n7242), .B(VbeatDelay_new_1_reg_326[20]), .C(
        VbeatDelay_new_1_reg_326[1]), .Y(n308) );
  NOR3X1 U76 ( .A(n7089), .B(VbeatDelay_new_1_reg_326[17]), .C(
        VbeatDelay_new_1_reg_326[16]), .Y(n307) );
  NAND3X1 U78 ( .A(n325), .B(n326), .C(n327), .Y(n305) );
  NOR3X1 U79 ( .A(n7611), .B(n7612), .C(n7610), .Y(n327) );
  NAND3X1 U81 ( .A(n10472), .B(n10474), .C(n10468), .Y(n329) );
  NAND3X1 U82 ( .A(n10531), .B(n10533), .C(n8018), .Y(n328) );
  NOR3X1 U84 ( .A(n6938), .B(VbeatDelay_new_1_reg_326[28]), .C(
        VbeatDelay_new_1_reg_326[27]), .Y(n326) );
  NOR3X1 U86 ( .A(n8022), .B(VbeatDelay_new_1_reg_326[24]), .C(
        VbeatDelay_new_1_reg_326[23]), .Y(n325) );
  AOI22X1 U89 ( .A(recentdatapoints_head_i[4]), .B(n367), .C(
        recentdatapoints_data_addr_reg_1533[4]), .D(ap_CS_fsm[1]), .Y(n347) );
  AOI22X1 U91 ( .A(p_tmp_i_reg_1556[4]), .B(n8397), .C(i_1_fu_620_p2[4]), .D(
        n9824), .Y(n345) );
  AOI22X1 U93 ( .A(recentdatapoints_head_i[3]), .B(n367), .C(
        recentdatapoints_data_addr_reg_1533[3]), .D(ap_CS_fsm[1]), .Y(n354) );
  AOI22X1 U95 ( .A(p_tmp_i_reg_1556[3]), .B(n8397), .C(i_1_fu_620_p2[3]), .D(
        n9824), .Y(n352) );
  AOI22X1 U97 ( .A(recentdatapoints_head_i[2]), .B(n367), .C(
        recentdatapoints_data_addr_reg_1533[2]), .D(ap_CS_fsm[1]), .Y(n357) );
  AOI22X1 U99 ( .A(p_tmp_i_reg_1556[2]), .B(n8397), .C(i_1_fu_620_p2[2]), .D(
        n9824), .Y(n355) );
  NAND3X1 U100 ( .A(n5451), .B(n5695), .C(n5860), .Y(
        recentdatapoints_data_address0[1]) );
  AOI22X1 U101 ( .A(recentdatapoints_head_i[1]), .B(n367), .C(
        recentdatapoints_data_addr_reg_1533[1]), .D(ap_CS_fsm[1]), .Y(n360) );
  AOI22X1 U103 ( .A(p_tmp_i_reg_1556[1]), .B(n8397), .C(i_1_fu_620_p2[1]), .D(
        n9824), .Y(n358) );
  NAND3X1 U104 ( .A(n5450), .B(n5694), .C(n5859), .Y(
        recentdatapoints_data_address0[0]) );
  AOI22X1 U105 ( .A(recentdatapoints_head_i[0]), .B(n367), .C(
        recentdatapoints_data_addr_reg_1533[0]), .D(ap_CS_fsm[1]), .Y(n363) );
  NOR3X1 U107 ( .A(n367), .B(i_fu_607_p2_31), .C(n8355), .Y(n349) );
  AOI22X1 U108 ( .A(p_tmp_i_reg_1556[0]), .B(n8397), .C(n9900), .D(n9824), .Y(
        n361) );
  NAND3X1 U110 ( .A(n364), .B(n8069), .C(i_fu_607_p2_31), .Y(n365) );
  AOI22X1 U113 ( .A(i_3_fu_835_p2[4]), .B(n371), .C(i_2_fu_823_p2[4]), .D(n372), .Y(n370) );
  AOI22X1 U114 ( .A(recentVBools_head_i[4]), .B(n373), .C(
        recentVBools_data_addr_reg_1573[4]), .D(n8981), .Y(n369) );
  AOI22X1 U116 ( .A(i_3_fu_835_p2[3]), .B(n371), .C(i_2_fu_823_p2[3]), .D(n372), .Y(n375) );
  AOI22X1 U117 ( .A(recentVBools_head_i[3]), .B(n373), .C(
        recentVBools_data_addr_reg_1573[3]), .D(n8981), .Y(n374) );
  AOI22X1 U119 ( .A(i_3_fu_835_p2[2]), .B(n371), .C(i_2_fu_823_p2[2]), .D(n372), .Y(n377) );
  AOI22X1 U120 ( .A(recentVBools_head_i[2]), .B(n373), .C(
        recentVBools_data_addr_reg_1573[2]), .D(n8981), .Y(n376) );
  AOI22X1 U122 ( .A(n9991), .B(n371), .C(i_2_fu_823_p2[1]), .D(n372), .Y(n379)
         );
  AOI22X1 U123 ( .A(recentVBools_head_i[1]), .B(n373), .C(
        recentVBools_data_addr_reg_1573[1]), .D(n8981), .Y(n378) );
  AOI22X1 U125 ( .A(i_3_fu_835_p2[0]), .B(n371), .C(i_3_fu_835_p2[0]), .D(n372), .Y(n381) );
  NOR3X1 U126 ( .A(n8981), .B(i_2_fu_823_p2[31]), .C(n373), .Y(n372) );
  NOR3X1 U127 ( .A(n373), .B(n8981), .C(n9965), .Y(n371) );
  AOI22X1 U129 ( .A(recentVBools_head_i[0]), .B(n373), .C(
        recentVBools_data_addr_reg_1573[0]), .D(n8981), .Y(n380) );
  AOI22X1 U131 ( .A(i_9_fu_1160_p2[4]), .B(n385), .C(i_8_fu_1148_p2[4]), .D(
        n386), .Y(n384) );
  AOI22X1 U132 ( .A(recentABools_head_i[4]), .B(n387), .C(
        recentABools_data_addr_reg_1689[4]), .D(ap_CS_fsm[9]), .Y(n383) );
  AOI22X1 U134 ( .A(i_9_fu_1160_p2[3]), .B(n385), .C(i_8_fu_1148_p2[3]), .D(
        n386), .Y(n389) );
  AOI22X1 U135 ( .A(recentABools_head_i[3]), .B(n387), .C(
        recentABools_data_addr_reg_1689[3]), .D(n9014), .Y(n388) );
  AOI22X1 U137 ( .A(i_9_fu_1160_p2[2]), .B(n385), .C(i_8_fu_1148_p2[2]), .D(
        n386), .Y(n391) );
  AOI22X1 U138 ( .A(recentABools_head_i[2]), .B(n387), .C(
        recentABools_data_addr_reg_1689[2]), .D(ap_CS_fsm[9]), .Y(n390) );
  AOI22X1 U140 ( .A(n10332), .B(n385), .C(i_8_fu_1148_p2[1]), .D(n386), .Y(
        n393) );
  AOI22X1 U141 ( .A(recentABools_head_i[1]), .B(n387), .C(
        recentABools_data_addr_reg_1689[1]), .D(ap_CS_fsm[9]), .Y(n392) );
  AOI22X1 U143 ( .A(i_9_fu_1160_p2[0]), .B(n385), .C(i_9_fu_1160_p2[0]), .D(
        n386), .Y(n395) );
  NOR3X1 U144 ( .A(n9014), .B(i_8_fu_1148_p2[31]), .C(n387), .Y(n386) );
  NOR3X1 U145 ( .A(n387), .B(n9014), .C(n10306), .Y(n385) );
  AOI22X1 U147 ( .A(recentABools_head_i[0]), .B(n387), .C(
        recentABools_data_addr_reg_1689[0]), .D(ap_CS_fsm[9]), .Y(n394) );
  OAI21X1 U148 ( .A(n397), .B(n8115), .C(n7380), .Y(p_cast_fu_688_p1_31) );
  OAI21X1 U150 ( .A(n397), .B(n7856), .C(n5198), .Y(p_cast_fu_688_p1[9]) );
  OAI21X1 U152 ( .A(n397), .B(n7436), .C(n5197), .Y(p_cast_fu_688_p1[8]) );
  OAI21X1 U154 ( .A(n397), .B(n7096), .C(n5196), .Y(p_cast_fu_688_p1[7]) );
  OAI21X1 U156 ( .A(n397), .B(n7435), .C(n5195), .Y(p_cast_fu_688_p1[6]) );
  OAI21X1 U158 ( .A(n397), .B(n7857), .C(n5194), .Y(p_cast_fu_688_p1[5]) );
  OAI21X1 U160 ( .A(n397), .B(n8101), .C(n5193), .Y(p_cast_fu_688_p1[4]) );
  OAI21X1 U162 ( .A(n397), .B(n7638), .C(n5192), .Y(p_cast_fu_688_p1[3]) );
  OAI21X1 U164 ( .A(n397), .B(n7261), .C(n5191), .Y(p_cast_fu_688_p1[2]) );
  OAI21X1 U166 ( .A(n397), .B(n6944), .C(n5190), .Y(p_cast_fu_688_p1[1]) );
  OAI21X1 U168 ( .A(n397), .B(n8115), .C(n5189), .Y(p_cast_fu_688_p1[15]) );
  OAI21X1 U170 ( .A(n397), .B(n6945), .C(n5188), .Y(p_cast_fu_688_p1[14]) );
  OAI21X1 U172 ( .A(n397), .B(n7639), .C(n5187), .Y(p_cast_fu_688_p1[13]) );
  OAI21X1 U174 ( .A(n397), .B(n8387), .C(n5186), .Y(p_cast_fu_688_p1[12]) );
  OAI21X1 U176 ( .A(n397), .B(n7262), .C(n5185), .Y(p_cast_fu_688_p1[11]) );
  OAI21X1 U178 ( .A(n397), .B(n7097), .C(n5184), .Y(p_cast_fu_688_p1[10]) );
  OAI21X1 U180 ( .A(n397), .B(n8390), .C(n7969), .Y(p_cast_fu_688_p1[0]) );
  NOR3X1 U183 ( .A(n8278), .B(n9542), .C(n9543), .Y(n432) );
  NOR3X1 U185 ( .A(n8020), .B(n9546), .C(n9547), .Y(n431) );
  OAI21X1 U187 ( .A(n439), .B(n8408), .C(n7381), .Y(p_1_cast_fu_1031_p1_31) );
  OAI21X1 U189 ( .A(n439), .B(n7263), .C(n5183), .Y(p_1_cast_fu_1031_p1[9]) );
  OAI21X1 U191 ( .A(n439), .B(n6811), .C(n5182), .Y(p_1_cast_fu_1031_p1[8]) );
  OAI21X1 U193 ( .A(n439), .B(n6164), .C(n5181), .Y(p_1_cast_fu_1031_p1[7]) );
  OAI21X1 U195 ( .A(n439), .B(n6571), .C(n5180), .Y(p_1_cast_fu_1031_p1[6]) );
  OAI21X1 U197 ( .A(n439), .B(n7437), .C(n5179), .Y(p_1_cast_fu_1031_p1[5]) );
  OAI21X1 U199 ( .A(n439), .B(n7640), .C(n5178), .Y(p_1_cast_fu_1031_p1[4]) );
  OAI21X1 U201 ( .A(n439), .B(n6946), .C(n5177), .Y(p_1_cast_fu_1031_p1[3]) );
  OAI21X1 U203 ( .A(n439), .B(n6458), .C(n5176), .Y(p_1_cast_fu_1031_p1[2]) );
  OAI21X1 U205 ( .A(n439), .B(n6093), .C(n5175), .Y(p_1_cast_fu_1031_p1[1]) );
  OAI21X1 U207 ( .A(n439), .B(n8408), .C(n5174), .Y(p_1_cast_fu_1031_p1[15])
         );
  OAI21X1 U209 ( .A(n439), .B(n6252), .C(n5173), .Y(p_1_cast_fu_1031_p1[14])
         );
  OAI21X1 U211 ( .A(n439), .B(n7098), .C(n5172), .Y(p_1_cast_fu_1031_p1[13])
         );
  OAI21X1 U213 ( .A(n439), .B(n7858), .C(n5171), .Y(p_1_cast_fu_1031_p1[12])
         );
  OAI21X1 U215 ( .A(n439), .B(n6686), .C(n5170), .Y(p_1_cast_fu_1031_p1[11])
         );
  OAI21X1 U217 ( .A(n439), .B(n6349), .C(n5169), .Y(p_1_cast_fu_1031_p1[10])
         );
  OAI21X1 U219 ( .A(n439), .B(n8107), .C(n7752), .Y(p_1_cast_fu_1031_p1[0]) );
  NOR3X1 U222 ( .A(n8279), .B(n9792), .C(n9491), .Y(n474) );
  NOR3X1 U224 ( .A(n8021), .B(n9494), .C(n9495), .Y(n473) );
  OAI21X1 U226 ( .A(n9040), .B(n4689), .C(n7720), .Y(n3257) );
  OAI21X1 U228 ( .A(n8974), .B(n10808), .C(n7936), .Y(n3258) );
  OAI21X1 U230 ( .A(ap_CS_fsm[12]), .B(n10809), .C(n7974), .Y(n3259) );
  OAI21X1 U233 ( .A(n8962), .B(n10808), .C(n8210), .Y(n3260) );
  OAI21X1 U236 ( .A(n8974), .B(n10807), .C(n8181), .Y(n3261) );
  OAI21X1 U238 ( .A(n8963), .B(n10807), .C(n7935), .Y(n3262) );
  OAI21X1 U241 ( .A(n8974), .B(n10806), .C(n7719), .Y(n3263) );
  OAI21X1 U243 ( .A(n8963), .B(n10806), .C(n8180), .Y(n3264) );
  OAI21X1 U246 ( .A(n8974), .B(n10805), .C(n7519), .Y(n3265) );
  OAI21X1 U248 ( .A(n8963), .B(n10805), .C(n7718), .Y(n3266) );
  OAI21X1 U251 ( .A(n8974), .B(n10804), .C(n7340), .Y(n3267) );
  OAI21X1 U253 ( .A(n8961), .B(n10804), .C(n7518), .Y(n3268) );
  OAI21X1 U256 ( .A(n8974), .B(n10803), .C(n7175), .Y(n3269) );
  OAI21X1 U258 ( .A(n8963), .B(n10803), .C(n7339), .Y(n3270) );
  OAI21X1 U261 ( .A(n8974), .B(n10802), .C(n7024), .Y(n3271) );
  OAI21X1 U263 ( .A(n8961), .B(n10802), .C(n7174), .Y(n3272) );
  OAI21X1 U266 ( .A(n8974), .B(n10801), .C(n6883), .Y(n3273) );
  OAI21X1 U268 ( .A(n8962), .B(n10801), .C(n7517), .Y(n3274) );
  OAI21X1 U271 ( .A(n8974), .B(n10800), .C(n7934), .Y(n3275) );
  OAI21X1 U273 ( .A(n8962), .B(n10800), .C(n7338), .Y(n3276) );
  OAI21X1 U276 ( .A(n8974), .B(n10799), .C(n8179), .Y(n3277) );
  OAI21X1 U278 ( .A(n8962), .B(n10799), .C(n7023), .Y(n3278) );
  OAI21X1 U281 ( .A(n8974), .B(n10798), .C(n7717), .Y(n3279) );
  OAI21X1 U283 ( .A(n8966), .B(n10798), .C(n6882), .Y(n3280) );
  OAI21X1 U286 ( .A(n8974), .B(n10797), .C(n7516), .Y(n3281) );
  OAI21X1 U288 ( .A(n8963), .B(n10797), .C(n6756), .Y(n3282) );
  OAI21X1 U291 ( .A(n8974), .B(n10796), .C(n7337), .Y(n3283) );
  OAI21X1 U293 ( .A(n8964), .B(n10796), .C(n6636), .Y(n3284) );
  OAI21X1 U296 ( .A(n8974), .B(n10795), .C(n7173), .Y(n3285) );
  OAI21X1 U298 ( .A(n8967), .B(n10795), .C(n6523), .Y(n3286) );
  OAI21X1 U301 ( .A(n8974), .B(n10794), .C(n6755), .Y(n3287) );
  OAI21X1 U303 ( .A(n8961), .B(n10794), .C(n6414), .Y(n3288) );
  OAI21X1 U306 ( .A(n8974), .B(n10793), .C(n6635), .Y(n3289) );
  OAI21X1 U308 ( .A(n8961), .B(n10793), .C(n6307), .Y(n3290) );
  OAI21X1 U311 ( .A(n8974), .B(n10792), .C(n6522), .Y(n3291) );
  OAI21X1 U313 ( .A(n8961), .B(n10792), .C(n6213), .Y(n3292) );
  OAI21X1 U316 ( .A(n8974), .B(n10791), .C(n6413), .Y(n3293) );
  OAI21X1 U318 ( .A(n8961), .B(n10791), .C(n6133), .Y(n3294) );
  OAI21X1 U321 ( .A(n8974), .B(n10790), .C(n6306), .Y(n3295) );
  OAI21X1 U323 ( .A(n8961), .B(n10790), .C(n6067), .Y(n3296) );
  OAI21X1 U326 ( .A(n8974), .B(n10789), .C(n6212), .Y(n3297) );
  OAI21X1 U328 ( .A(n8965), .B(n10789), .C(n5168), .Y(n3298) );
  OAI21X1 U331 ( .A(n8974), .B(n10788), .C(n6132), .Y(n3299) );
  OAI21X1 U333 ( .A(n8658), .B(n10788), .C(n5167), .Y(n3300) );
  OAI21X1 U336 ( .A(n8974), .B(n10787), .C(n6066), .Y(n3301) );
  OAI21X1 U338 ( .A(n8962), .B(n10787), .C(n7933), .Y(n3302) );
  OAI21X1 U341 ( .A(n8974), .B(n10786), .C(n5166), .Y(n3303) );
  OAI21X1 U343 ( .A(n8962), .B(n10786), .C(n7172), .Y(n3304) );
  OAI21X1 U346 ( .A(n8974), .B(n10785), .C(n8178), .Y(n3305) );
  OAI21X1 U348 ( .A(n8961), .B(n10785), .C(n7515), .Y(n3306) );
  OAI21X1 U351 ( .A(n8974), .B(n10784), .C(n7932), .Y(n3307) );
  OAI21X1 U353 ( .A(n8963), .B(n10784), .C(n7336), .Y(n3308) );
  OAI21X1 U356 ( .A(n8974), .B(n10783), .C(n7716), .Y(n3309) );
  OAI21X1 U358 ( .A(n8967), .B(n10783), .C(n7022), .Y(n3310) );
  OAI21X1 U361 ( .A(n8974), .B(n10782), .C(n7514), .Y(n3311) );
  OAI21X1 U363 ( .A(n8964), .B(n10782), .C(n6881), .Y(n3312) );
  OAI21X1 U366 ( .A(n8974), .B(n10781), .C(n7335), .Y(n3313) );
  OAI21X1 U368 ( .A(n8966), .B(n10781), .C(n6754), .Y(n3314) );
  OAI21X1 U371 ( .A(n8974), .B(n10780), .C(n7171), .Y(n3315) );
  OAI21X1 U373 ( .A(n8962), .B(n10780), .C(n6634), .Y(n3316) );
  OAI21X1 U376 ( .A(n8974), .B(n10779), .C(n7021), .Y(n3317) );
  OAI21X1 U378 ( .A(n8961), .B(n10779), .C(n6521), .Y(n3318) );
  OAI21X1 U381 ( .A(n8974), .B(n10778), .C(n6880), .Y(n3319) );
  OAI21X1 U383 ( .A(n8961), .B(n10778), .C(n6412), .Y(n3320) );
  OAI21X1 U386 ( .A(n8961), .B(n10777), .C(n5165), .Y(n3321) );
  OAI21X1 U388 ( .A(n8974), .B(n10777), .C(n6753), .Y(n3322) );
  OAI21X1 U392 ( .A(n8973), .B(n10774), .C(n6752), .Y(n3323) );
  OAI21X1 U394 ( .A(ap_CS_fsm[12]), .B(n10775), .C(n7757), .Y(n3324) );
  OAI21X1 U397 ( .A(n8961), .B(n10774), .C(n7751), .Y(n3325) );
  OAI21X1 U400 ( .A(n8973), .B(n10773), .C(n6633), .Y(n3326) );
  OAI21X1 U402 ( .A(n8961), .B(n10773), .C(n5164), .Y(n3327) );
  OAI21X1 U405 ( .A(n8973), .B(n10772), .C(n6520), .Y(n3328) );
  OAI21X1 U407 ( .A(n8961), .B(n10772), .C(n5163), .Y(n3329) );
  OAI21X1 U410 ( .A(n8973), .B(n10771), .C(n6411), .Y(n3330) );
  OAI21X1 U412 ( .A(n8961), .B(n10771), .C(n5162), .Y(n3331) );
  OAI21X1 U415 ( .A(n8973), .B(n10770), .C(n6305), .Y(n3332) );
  OAI21X1 U417 ( .A(n8961), .B(n10770), .C(n5161), .Y(n3333) );
  OAI21X1 U420 ( .A(n8973), .B(n10769), .C(n6211), .Y(n3334) );
  OAI21X1 U422 ( .A(n8961), .B(n10769), .C(n8177), .Y(n3335) );
  OAI21X1 U425 ( .A(n8973), .B(n10768), .C(n6131), .Y(n3336) );
  OAI21X1 U427 ( .A(n8963), .B(n10768), .C(n7931), .Y(n3337) );
  OAI21X1 U430 ( .A(n8973), .B(n10767), .C(n6065), .Y(n3338) );
  OAI21X1 U432 ( .A(n8658), .B(n10767), .C(n7715), .Y(n3339) );
  OAI21X1 U435 ( .A(n8973), .B(n10766), .C(n5160), .Y(n3340) );
  OAI21X1 U437 ( .A(n8966), .B(n10766), .C(n7513), .Y(n3341) );
  OAI21X1 U440 ( .A(n8973), .B(n10765), .C(n8176), .Y(n3342) );
  OAI21X1 U442 ( .A(n8965), .B(n10765), .C(n7334), .Y(n3343) );
  OAI21X1 U445 ( .A(n8973), .B(n10764), .C(n7930), .Y(n3344) );
  OAI21X1 U447 ( .A(n8962), .B(n10764), .C(n7170), .Y(n3345) );
  OAI21X1 U450 ( .A(n8973), .B(n10763), .C(n7714), .Y(n3346) );
  OAI21X1 U452 ( .A(n8961), .B(n10763), .C(n7020), .Y(n3347) );
  OAI21X1 U455 ( .A(n8973), .B(n10762), .C(n7512), .Y(n3348) );
  OAI21X1 U457 ( .A(n8658), .B(n10762), .C(n6304), .Y(n3349) );
  OAI21X1 U460 ( .A(n8973), .B(n10761), .C(n7333), .Y(n3350) );
  OAI21X1 U462 ( .A(n8967), .B(n10761), .C(n6210), .Y(n3351) );
  OAI21X1 U465 ( .A(n8973), .B(n10760), .C(n7169), .Y(n3352) );
  OAI21X1 U467 ( .A(n8962), .B(n10760), .C(n6879), .Y(n3353) );
  OAI21X1 U470 ( .A(n8973), .B(n10759), .C(n7019), .Y(n3354) );
  OAI21X1 U472 ( .A(n8962), .B(n10759), .C(n6751), .Y(n3355) );
  OAI21X1 U475 ( .A(n8973), .B(n10758), .C(n6878), .Y(n3356) );
  OAI21X1 U477 ( .A(n8962), .B(n10758), .C(n6632), .Y(n3357) );
  OAI21X1 U480 ( .A(n8973), .B(n10757), .C(n6750), .Y(n3358) );
  OAI21X1 U482 ( .A(n8962), .B(n10757), .C(n6519), .Y(n3359) );
  OAI21X1 U485 ( .A(n8973), .B(n10756), .C(n6631), .Y(n3360) );
  OAI21X1 U487 ( .A(n8962), .B(n10756), .C(n6410), .Y(n3361) );
  OAI21X1 U490 ( .A(n8973), .B(n10755), .C(n6518), .Y(n3362) );
  OAI21X1 U492 ( .A(n8962), .B(n10755), .C(n6130), .Y(n3363) );
  OAI21X1 U495 ( .A(n8973), .B(n10754), .C(n6409), .Y(n3364) );
  OAI21X1 U497 ( .A(n8962), .B(n10754), .C(n6064), .Y(n3365) );
  OAI21X1 U500 ( .A(n8973), .B(n10753), .C(n6303), .Y(n3366) );
  OAI21X1 U502 ( .A(n8962), .B(n10753), .C(n5159), .Y(n3367) );
  OAI21X1 U505 ( .A(n8973), .B(n10752), .C(n6209), .Y(n3368) );
  OAI21X1 U507 ( .A(n8962), .B(n10752), .C(n5158), .Y(n3369) );
  OAI21X1 U510 ( .A(n8973), .B(n10751), .C(n6129), .Y(n3370) );
  OAI21X1 U512 ( .A(n8967), .B(n10751), .C(n8175), .Y(n3371) );
  OAI21X1 U515 ( .A(n8973), .B(n10750), .C(n6063), .Y(n3372) );
  OAI21X1 U517 ( .A(n8658), .B(n10750), .C(n7929), .Y(n3373) );
  OAI21X1 U520 ( .A(n8973), .B(n10749), .C(n5157), .Y(n3374) );
  OAI21X1 U522 ( .A(n8961), .B(n10749), .C(n7713), .Y(n3375) );
  OAI21X1 U525 ( .A(n8973), .B(n10748), .C(n8174), .Y(n3376) );
  OAI21X1 U527 ( .A(n8967), .B(n10748), .C(n6302), .Y(n3377) );
  OAI21X1 U530 ( .A(n8973), .B(n10747), .C(n7928), .Y(n3378) );
  OAI21X1 U532 ( .A(n8658), .B(n10747), .C(n7018), .Y(n3379) );
  OAI21X1 U535 ( .A(n8973), .B(n10746), .C(n7712), .Y(n3380) );
  OAI21X1 U537 ( .A(n8967), .B(n10746), .C(n6877), .Y(n3381) );
  OAI21X1 U540 ( .A(n8973), .B(n10745), .C(n7511), .Y(n3382) );
  OAI21X1 U542 ( .A(n8963), .B(n10745), .C(n7168), .Y(n3383) );
  OAI21X1 U545 ( .A(n8973), .B(n10744), .C(n7332), .Y(n3384) );
  OAI21X1 U547 ( .A(n8965), .B(n10744), .C(n6749), .Y(n3385) );
  OAI21X1 U550 ( .A(n8963), .B(n10743), .C(n6630), .Y(n3386) );
  OAI21X1 U552 ( .A(n8973), .B(n10743), .C(n7167), .Y(n3387) );
  OAI21X1 U556 ( .A(n10670), .B(n10741), .C(n7017), .Y(n3388) );
  OAI21X1 U559 ( .A(n8989), .B(n10740), .C(n7927), .Y(n3389) );
  OAI21X1 U561 ( .A(n10670), .B(n10739), .C(n6876), .Y(n3390) );
  OAI21X1 U564 ( .A(n8987), .B(n10738), .C(n7711), .Y(n3391) );
  OAI21X1 U566 ( .A(n8896), .B(n10737), .C(n6629), .Y(n3392) );
  OAI21X1 U569 ( .A(n8987), .B(n10736), .C(n8171), .Y(n3393) );
  OAI21X1 U571 ( .A(n10670), .B(n10735), .C(n6517), .Y(n3394) );
  OAI21X1 U574 ( .A(n8987), .B(n10734), .C(n7925), .Y(n3395) );
  OAI21X1 U576 ( .A(n8896), .B(n10733), .C(n6408), .Y(n3396) );
  OAI21X1 U579 ( .A(n8987), .B(n10732), .C(n7331), .Y(n3397) );
  OAI21X1 U581 ( .A(n8896), .B(n10731), .C(n6301), .Y(n3398) );
  OAI21X1 U584 ( .A(n8987), .B(n10730), .C(n7509), .Y(n3399) );
  OAI21X1 U586 ( .A(n8896), .B(n10729), .C(n6208), .Y(n3400) );
  OAI21X1 U589 ( .A(n8987), .B(n10728), .C(n7016), .Y(n3401) );
  OAI21X1 U591 ( .A(n10670), .B(n10727), .C(n8170), .Y(n3402) );
  OAI21X1 U594 ( .A(n8987), .B(n10726), .C(n7165), .Y(n3403) );
  OAI21X1 U596 ( .A(n10670), .B(n10725), .C(n7508), .Y(n3404) );
  OAI21X1 U599 ( .A(n8988), .B(n10724), .C(n7709), .Y(n3405) );
  OAI21X1 U601 ( .A(n8896), .B(n10723), .C(n7708), .Y(n3406) );
  OAI21X1 U604 ( .A(n8988), .B(n10722), .C(n6874), .Y(n3407) );
  OAI21X1 U606 ( .A(n10670), .B(n10721), .C(n6128), .Y(n3408) );
  OAI21X1 U609 ( .A(n8988), .B(n10720), .C(n6747), .Y(n3409) );
  OAI21X1 U611 ( .A(n8896), .B(n10719), .C(n7329), .Y(n3410) );
  OAI21X1 U614 ( .A(n8988), .B(n10718), .C(n6627), .Y(n3411) );
  OAI21X1 U616 ( .A(n10670), .B(n10717), .C(n7164), .Y(n3412) );
  OAI21X1 U619 ( .A(n8988), .B(n10716), .C(n6515), .Y(n3413) );
  OAI21X1 U621 ( .A(n10670), .B(n10715), .C(n6062), .Y(n3414) );
  OAI21X1 U624 ( .A(n8988), .B(n10714), .C(n6406), .Y(n3415) );
  OAI21X1 U626 ( .A(n10670), .B(n10713), .C(n6873), .Y(n3416) );
  OAI21X1 U629 ( .A(n8988), .B(n10712), .C(n6300), .Y(n3417) );
  OAI21X1 U631 ( .A(n10670), .B(n10711), .C(n6746), .Y(n3418) );
  OAI21X1 U634 ( .A(n8988), .B(n10710), .C(n6207), .Y(n3419) );
  OAI21X1 U636 ( .A(n10670), .B(n10709), .C(n6626), .Y(n3420) );
  OAI21X1 U639 ( .A(n8988), .B(n10708), .C(n6127), .Y(n3421) );
  OAI21X1 U641 ( .A(n10670), .B(n10707), .C(n6405), .Y(n3422) );
  OAI21X1 U644 ( .A(n8988), .B(n10706), .C(n6061), .Y(n3423) );
  OAI21X1 U646 ( .A(n10670), .B(n10705), .C(n6299), .Y(n3424) );
  OAI21X1 U649 ( .A(n8989), .B(n10704), .C(n5156), .Y(n3425) );
  OAI21X1 U651 ( .A(n8896), .B(n10703), .C(n5155), .Y(n3426) );
  OAI21X1 U654 ( .A(n8989), .B(n10702), .C(n5154), .Y(n3427) );
  OAI21X1 U656 ( .A(n10670), .B(n10701), .C(n7014), .Y(n3428) );
  OAI21X1 U659 ( .A(n8989), .B(n10700), .C(n5153), .Y(n3429) );
  OAI21X1 U661 ( .A(n10670), .B(n10699), .C(n6205), .Y(n3430) );
  OAI21X1 U664 ( .A(n8989), .B(n10698), .C(n7706), .Y(n3431) );
  OAI21X1 U666 ( .A(n8896), .B(n10697), .C(n6514), .Y(n3432) );
  OAI21X1 U669 ( .A(n8989), .B(n10696), .C(n7506), .Y(n3433) );
  OAI21X1 U671 ( .A(n8896), .B(n10695), .C(n6125), .Y(n3434) );
  OAI21X1 U674 ( .A(n8989), .B(n10694), .C(n7327), .Y(n3435) );
  OAI21X1 U676 ( .A(n10670), .B(n10693), .C(n6060), .Y(n3436) );
  OAI21X1 U679 ( .A(n8989), .B(n10692), .C(n7162), .Y(n3437) );
  OAI21X1 U681 ( .A(n8896), .B(n10691), .C(n8168), .Y(n3438) );
  OAI21X1 U684 ( .A(n8990), .B(n10690), .C(n7012), .Y(n3439) );
  OAI21X1 U686 ( .A(n10670), .B(n10689), .C(n7922), .Y(n3440) );
  OAI21X1 U689 ( .A(n8989), .B(n10687), .C(n6871), .Y(n3441) );
  OAI21X1 U691 ( .A(n8896), .B(n10686), .C(n5152), .Y(n3442) );
  OAI21X1 U694 ( .A(n8990), .B(n10684), .C(n7921), .Y(n3443) );
  OAI21X1 U696 ( .A(n10670), .B(n10683), .C(n7504), .Y(n3444) );
  OAI21X1 U699 ( .A(n8990), .B(n10682), .C(n6744), .Y(n3445) );
  OAI21X1 U701 ( .A(n10670), .B(n10681), .C(n7161), .Y(n3446) );
  OAI21X1 U704 ( .A(n8990), .B(n10680), .C(n8167), .Y(n3447) );
  OAI21X1 U706 ( .A(n8896), .B(n10679), .C(n6743), .Y(n3448) );
  OAI21X1 U709 ( .A(n8991), .B(n10678), .C(n6513), .Y(n3449) );
  OAI21X1 U711 ( .A(n8990), .B(n10672), .C(n6624), .Y(n3450) );
  OAI21X1 U713 ( .A(n10670), .B(n10677), .C(n5151), .Y(n3451) );
  AOI22X1 U716 ( .A(n794), .B(n795), .C(n10534), .D(n10668), .Y(n3452) );
  NOR3X1 U718 ( .A(n7237), .B(n7608), .C(n8045), .Y(n795) );
  NAND3X1 U719 ( .A(n10657), .B(n10658), .C(n8046), .Y(n800) );
  NAND3X1 U721 ( .A(n10661), .B(n10662), .C(n7609), .Y(n799) );
  NOR3X1 U724 ( .A(n7238), .B(CircularBuffer_len_write_assig_2_reg_1729[6]), 
        .C(CircularBuffer_len_write_assig_2_reg_1729[5]), .Y(n808) );
  NAND3X1 U725 ( .A(n10642), .B(n10643), .C(n10641), .Y(n809) );
  NOR3X1 U726 ( .A(n8281), .B(CircularBuffer_len_write_assig_2_reg_1729[31]), 
        .C(CircularBuffer_len_write_assig_2_reg_1729[30]), .Y(n807) );
  NOR3X1 U728 ( .A(n7413), .B(n7808), .C(n8288), .Y(n794) );
  NAND3X1 U729 ( .A(n10650), .B(n10651), .C(n8289), .Y(n818) );
  NAND3X1 U731 ( .A(n10635), .B(n10654), .C(n7809), .Y(n817) );
  NOR3X1 U734 ( .A(n7414), .B(CircularBuffer_len_write_assig_2_reg_1729[13]), 
        .C(CircularBuffer_len_write_assig_2_reg_1729[12]), .Y(n826) );
  NOR3X1 U736 ( .A(n8273), .B(CircularBuffer_len_write_assig_2_reg_1729[11]), 
        .C(CircularBuffer_len_write_assig_2_reg_1729[10]), .Y(n825) );
  OAI21X1 U738 ( .A(n11047), .B(n833), .C(n7079), .Y(n3453) );
  OAI21X1 U740 ( .A(n7080), .B(n7234), .C(ap_CS_fsm[11]), .Y(n833) );
  NAND3X1 U741 ( .A(n838), .B(n839), .C(n840), .Y(n837) );
  NOR3X1 U742 ( .A(n8276), .B(n7803), .C(n8039), .Y(n840) );
  NAND3X1 U745 ( .A(n10593), .B(n10594), .C(n8277), .Y(n841) );
  NOR3X1 U747 ( .A(n7601), .B(CircularBuffer_len_read_assign_3_reg_1711[14]), 
        .C(CircularBuffer_len_read_assign_3_reg_1711[13]), .Y(n839) );
  NOR3X1 U749 ( .A(n7410), .B(CircularBuffer_len_read_assign_3_reg_1711[10]), 
        .C(CircularBuffer_len_write_assig_3_fu_1249_p2[0]), .Y(n838) );
  NAND3X1 U751 ( .A(n857), .B(n858), .C(n859), .Y(n836) );
  NOR3X1 U752 ( .A(n7812), .B(n7810), .C(n7811), .Y(n859) );
  NAND3X1 U755 ( .A(n10579), .B(n10580), .C(n8252), .Y(n860) );
  NOR3X1 U757 ( .A(n8019), .B(CircularBuffer_len_read_assign_3_reg_1711[29]), 
        .C(CircularBuffer_len_read_assign_3_reg_1711[28]), .Y(n858) );
  NOR3X1 U759 ( .A(n8271), .B(CircularBuffer_len_read_assign_3_reg_1711[25]), 
        .C(CircularBuffer_len_read_assign_3_reg_1711[24]), .Y(n857) );
  OAI21X1 U761 ( .A(n11047), .B(n10242), .C(n8165), .Y(n3454) );
  OAI21X1 U764 ( .A(n8891), .B(n10665), .C(n5150), .Y(n3455) );
  OAI21X1 U767 ( .A(n8891), .B(n10664), .C(n7920), .Y(n3456) );
  OAI21X1 U770 ( .A(n8891), .B(n10663), .C(n5149), .Y(n3457) );
  OAI21X1 U773 ( .A(n970), .B(n10662), .C(n5148), .Y(n3458) );
  OAI21X1 U776 ( .A(n8891), .B(n10661), .C(n5147), .Y(n3459) );
  OAI21X1 U779 ( .A(n970), .B(n10660), .C(n5146), .Y(n3460) );
  OAI21X1 U782 ( .A(n970), .B(n10659), .C(n5145), .Y(n3461) );
  OAI21X1 U785 ( .A(n8891), .B(n10658), .C(n5144), .Y(n3462) );
  OAI21X1 U788 ( .A(n970), .B(n10657), .C(n7503), .Y(n3463) );
  OAI21X1 U791 ( .A(n8891), .B(n10656), .C(n5143), .Y(n3464) );
  OAI21X1 U794 ( .A(n970), .B(n10655), .C(n5142), .Y(n3465) );
  OAI21X1 U797 ( .A(n970), .B(n10654), .C(n5141), .Y(n3466) );
  OAI21X1 U800 ( .A(n970), .B(n10653), .C(n5140), .Y(n3467) );
  OAI21X1 U803 ( .A(n8891), .B(n10652), .C(n5139), .Y(n3468) );
  OAI21X1 U806 ( .A(n970), .B(n10651), .C(n5138), .Y(n3469) );
  OAI21X1 U809 ( .A(n8891), .B(n10650), .C(n5137), .Y(n3470) );
  OAI21X1 U812 ( .A(n8891), .B(n10649), .C(n7011), .Y(n3471) );
  OAI21X1 U815 ( .A(n970), .B(n10648), .C(n6870), .Y(n3472) );
  OAI21X1 U818 ( .A(n970), .B(n10647), .C(n5136), .Y(n3473) );
  OAI21X1 U821 ( .A(n8891), .B(n10646), .C(n5135), .Y(n3474) );
  OAI21X1 U824 ( .A(n970), .B(n10645), .C(n7559), .Y(n3475) );
  OAI21X1 U827 ( .A(n970), .B(n10644), .C(n7218), .Y(n3476) );
  OAI21X1 U830 ( .A(n970), .B(n10643), .C(n7325), .Y(n3477) );
  OAI21X1 U833 ( .A(n970), .B(n10642), .C(n7703), .Y(n3478) );
  OAI21X1 U836 ( .A(n8891), .B(n10641), .C(n6742), .Y(n3479) );
  OAI21X1 U839 ( .A(n970), .B(n10640), .C(n5134), .Y(n3480) );
  OAI21X1 U842 ( .A(n970), .B(n10639), .C(n7010), .Y(n3481) );
  OAI21X1 U845 ( .A(n970), .B(n10638), .C(n6869), .Y(n3482) );
  OAI21X1 U848 ( .A(n8891), .B(n10637), .C(n6741), .Y(n3483) );
  OAI21X1 U851 ( .A(n8891), .B(n10636), .C(n6623), .Y(n3484) );
  OAI21X1 U854 ( .A(n970), .B(n10635), .C(n6511), .Y(n3485) );
  OAI21X1 U857 ( .A(n970), .B(n10634), .C(n6404), .Y(n3486) );
  OAI21X1 U860 ( .A(ap_CS_fsm[9]), .B(n10604), .C(n7916), .Y(n3487) );
  OAI21X1 U863 ( .A(n9015), .B(n10603), .C(n7700), .Y(n3488) );
  OAI21X1 U866 ( .A(n9016), .B(n10602), .C(n5133), .Y(n3489) );
  OAI21X1 U869 ( .A(ap_CS_fsm[9]), .B(n10601), .C(n5132), .Y(n3490) );
  OAI21X1 U872 ( .A(n9015), .B(n10600), .C(n7155), .Y(n3491) );
  OAI21X1 U875 ( .A(n9014), .B(n10599), .C(n5131), .Y(n3492) );
  OAI21X1 U878 ( .A(ap_CS_fsm[9]), .B(n10598), .C(n5130), .Y(n3493) );
  OAI21X1 U881 ( .A(n9014), .B(n10597), .C(n5129), .Y(n3494) );
  OAI21X1 U884 ( .A(n9015), .B(n10596), .C(n7318), .Y(n3495) );
  OAI21X1 U887 ( .A(n9015), .B(n10595), .C(n6865), .Y(n3496) );
  OAI21X1 U890 ( .A(n9015), .B(n10594), .C(n5128), .Y(n3497) );
  OAI21X1 U893 ( .A(n9015), .B(n10593), .C(n5127), .Y(n3498) );
  OAI21X1 U896 ( .A(n9015), .B(n10592), .C(n5126), .Y(n3499) );
  OAI21X1 U899 ( .A(n9015), .B(n10591), .C(n5125), .Y(n3500) );
  OAI21X1 U902 ( .A(n9015), .B(n10590), .C(n5124), .Y(n3501) );
  OAI21X1 U905 ( .A(n9015), .B(n10589), .C(n5123), .Y(n3502) );
  OAI21X1 U908 ( .A(n9016), .B(n10588), .C(n7154), .Y(n3503) );
  OAI21X1 U911 ( .A(n9016), .B(n10587), .C(n7496), .Y(n3504) );
  OAI21X1 U914 ( .A(n9016), .B(n10586), .C(n5122), .Y(n3505) );
  OAI21X1 U917 ( .A(n9016), .B(n10585), .C(n5121), .Y(n3506) );
  OAI21X1 U920 ( .A(n9015), .B(n10584), .C(n7005), .Y(n3507) );
  OAI21X1 U923 ( .A(n9017), .B(n10583), .C(n7317), .Y(n3508) );
  OAI21X1 U926 ( .A(n9017), .B(n10582), .C(n6737), .Y(n3509) );
  OAI21X1 U929 ( .A(n9017), .B(n10581), .C(n6507), .Y(n3510) );
  OAI21X1 U932 ( .A(n9016), .B(n10580), .C(n6400), .Y(n3511) );
  OAI21X1 U935 ( .A(n9017), .B(n10579), .C(n5120), .Y(n3512) );
  OAI21X1 U938 ( .A(n9015), .B(n10578), .C(n5119), .Y(n3513) );
  OAI21X1 U941 ( .A(n9016), .B(n10577), .C(n8163), .Y(n3514) );
  OAI21X1 U944 ( .A(n9016), .B(n10576), .C(n7915), .Y(n3515) );
  OAI21X1 U947 ( .A(n9016), .B(n10575), .C(n7699), .Y(n3516) );
  OAI21X1 U950 ( .A(n9016), .B(n10574), .C(n7004), .Y(n3517) );
  OAI21X1 U953 ( .A(n9017), .B(n10542), .C(n8892), .Y(n3518) );
  OAI21X1 U955 ( .A(n9017), .B(n10541), .C(n6291), .Y(n3519) );
  OAI21X1 U958 ( .A(n9021), .B(n10533), .C(n8161), .Y(n3520) );
  OAI21X1 U961 ( .A(n8990), .B(n10532), .C(n6395), .Y(n3521) );
  OAI21X1 U963 ( .A(n9027), .B(n10531), .C(n8160), .Y(n3522) );
  OAI21X1 U966 ( .A(n8990), .B(n10528), .C(n6290), .Y(n3523) );
  OAI21X1 U968 ( .A(n9027), .B(n10527), .C(n7911), .Y(n3524) );
  OAI21X1 U971 ( .A(n8990), .B(n10526), .C(n6199), .Y(n3525) );
  OAI21X1 U973 ( .A(n9027), .B(n10525), .C(n7694), .Y(n3526) );
  OAI21X1 U976 ( .A(n8990), .B(n10524), .C(n6123), .Y(n3527) );
  OAI21X1 U978 ( .A(n9027), .B(n10523), .C(n7491), .Y(n3528) );
  OAI21X1 U981 ( .A(n8991), .B(n10522), .C(n6058), .Y(n3529) );
  OAI21X1 U983 ( .A(n9027), .B(n10521), .C(n7311), .Y(n3530) );
  OAI21X1 U986 ( .A(n8989), .B(n10518), .C(n5118), .Y(n3531) );
  OAI21X1 U988 ( .A(n9026), .B(n10517), .C(n8158), .Y(n3532) );
  OAI21X1 U991 ( .A(n8986), .B(n10516), .C(n5117), .Y(n3533) );
  OAI21X1 U993 ( .A(n9026), .B(n10515), .C(n7909), .Y(n3534) );
  OAI21X1 U996 ( .A(n8986), .B(n10513), .C(n5116), .Y(n3535) );
  OAI21X1 U998 ( .A(n9026), .B(n10512), .C(n7693), .Y(n3536) );
  OAI21X1 U1001 ( .A(n8986), .B(n10511), .C(n8157), .Y(n3537) );
  OAI21X1 U1003 ( .A(n9026), .B(n10510), .C(n7490), .Y(n3538) );
  OAI21X1 U1006 ( .A(n8986), .B(n10507), .C(n7908), .Y(n3539) );
  OAI21X1 U1008 ( .A(n9026), .B(n10506), .C(n7310), .Y(n3540) );
  OAI21X1 U1011 ( .A(n8986), .B(n10505), .C(n7692), .Y(n3541) );
  OAI21X1 U1013 ( .A(n9026), .B(n10504), .C(n6997), .Y(n3542) );
  OAI21X1 U1016 ( .A(n8986), .B(n10502), .C(n7489), .Y(n3543) );
  OAI21X1 U1018 ( .A(n9026), .B(n10501), .C(n7146), .Y(n3544) );
  OAI21X1 U1021 ( .A(n8986), .B(n10500), .C(n7309), .Y(n3545) );
  OAI21X1 U1023 ( .A(n9026), .B(n10499), .C(n6857), .Y(n3546) );
  OAI21X1 U1026 ( .A(n8986), .B(n10496), .C(n7145), .Y(n3547) );
  OAI21X1 U1028 ( .A(n9026), .B(n10495), .C(n6729), .Y(n3548) );
  OAI21X1 U1031 ( .A(n8986), .B(n10494), .C(n6996), .Y(n3549) );
  OAI21X1 U1033 ( .A(n9026), .B(n10493), .C(n6612), .Y(n3550) );
  OAI21X1 U1036 ( .A(n8985), .B(n10492), .C(n6856), .Y(n3551) );
  OAI21X1 U1038 ( .A(n9026), .B(n10491), .C(n6500), .Y(n3552) );
  OAI21X1 U1041 ( .A(n8985), .B(n10490), .C(n6728), .Y(n3553) );
  OAI21X1 U1043 ( .A(n9026), .B(n10489), .C(n6393), .Y(n3554) );
  OAI21X1 U1046 ( .A(n8985), .B(n10486), .C(n6611), .Y(n3555) );
  OAI21X1 U1048 ( .A(n9025), .B(n10485), .C(n8155), .Y(n3556) );
  OAI21X1 U1051 ( .A(n8985), .B(n10484), .C(n6499), .Y(n3557) );
  OAI21X1 U1053 ( .A(n9025), .B(n10483), .C(n7307), .Y(n3558) );
  OAI21X1 U1056 ( .A(n8985), .B(n10481), .C(n6392), .Y(n3559) );
  OAI21X1 U1058 ( .A(n9025), .B(n10480), .C(n6994), .Y(n3560) );
  OAI21X1 U1061 ( .A(n8985), .B(n10479), .C(n6289), .Y(n3561) );
  OAI21X1 U1063 ( .A(n9025), .B(n10478), .C(n6610), .Y(n3562) );
  OAI21X1 U1066 ( .A(n8985), .B(n10475), .C(n6198), .Y(n3563) );
  OAI21X1 U1068 ( .A(n9025), .B(n10474), .C(n7143), .Y(n3564) );
  OAI21X1 U1071 ( .A(n8985), .B(n10473), .C(n6122), .Y(n3565) );
  OAI21X1 U1073 ( .A(n9025), .B(n10472), .C(n7906), .Y(n3566) );
  OAI21X1 U1076 ( .A(n8985), .B(n10469), .C(n6057), .Y(n3567) );
  OAI21X1 U1078 ( .A(n9025), .B(n10468), .C(n7690), .Y(n3568) );
  OAI21X1 U1081 ( .A(n8984), .B(n10467), .C(n5115), .Y(n3569) );
  OAI21X1 U1083 ( .A(n9025), .B(n10466), .C(n6854), .Y(n3570) );
  OAI21X1 U1086 ( .A(n8984), .B(n10464), .C(n5114), .Y(n3571) );
  OAI21X1 U1088 ( .A(n9025), .B(n10463), .C(n6726), .Y(n3572) );
  OAI21X1 U1091 ( .A(n8984), .B(n10462), .C(n5113), .Y(n3573) );
  OAI21X1 U1093 ( .A(n9025), .B(n10461), .C(n7486), .Y(n3574) );
  OAI21X1 U1096 ( .A(n8984), .B(n10460), .C(n8153), .Y(n3575) );
  OAI21X1 U1098 ( .A(n8984), .B(n10458), .C(n7904), .Y(n3576) );
  OAI21X1 U1100 ( .A(n9025), .B(n10457), .C(n6497), .Y(n3577) );
  OAI21X1 U1103 ( .A(n8984), .B(n10455), .C(n7688), .Y(n3578) );
  OAI21X1 U1105 ( .A(n9025), .B(n10454), .C(n6390), .Y(n3579) );
  OAI21X1 U1108 ( .A(n8984), .B(n10453), .C(n7485), .Y(n3580) );
  OAI21X1 U1110 ( .A(n9024), .B(n10451), .C(n6992), .Y(n3581) );
  OAI21X1 U1113 ( .A(n8984), .B(n10450), .C(n7305), .Y(n3582) );
  OAI21X1 U1115 ( .A(n9024), .B(n10459), .C(n6608), .Y(n3583) );
  OAI21X1 U1118 ( .A(n9024), .B(n10449), .C(n7304), .Y(n3584) );
  OAI21X1 U1121 ( .A(n8984), .B(n10448), .C(n7141), .Y(n3585) );
  OAI21X1 U1123 ( .A(n9024), .B(n10447), .C(n7140), .Y(n3586) );
  OAI21X1 U1126 ( .A(n8984), .B(n10444), .C(n6991), .Y(n3587) );
  OAI21X1 U1128 ( .A(n9024), .B(n10443), .C(n6852), .Y(n3588) );
  OAI21X1 U1131 ( .A(n8983), .B(n10442), .C(n6851), .Y(n3589) );
  OAI21X1 U1133 ( .A(n9024), .B(n10441), .C(n6725), .Y(n3590) );
  OAI21X1 U1136 ( .A(n8983), .B(n10440), .C(n6724), .Y(n3591) );
  OAI21X1 U1138 ( .A(n9024), .B(n10439), .C(n6496), .Y(n3592) );
  OAI21X1 U1141 ( .A(n8983), .B(n10438), .C(n6607), .Y(n3593) );
  OAI21X1 U1143 ( .A(n9024), .B(n10437), .C(n6389), .Y(n3594) );
  OAI21X1 U1146 ( .A(n8983), .B(n10434), .C(n6495), .Y(n3595) );
  OAI21X1 U1148 ( .A(n9024), .B(n10433), .C(n6288), .Y(n3596) );
  OAI21X1 U1151 ( .A(n8983), .B(n10432), .C(n6388), .Y(n3597) );
  OAI21X1 U1153 ( .A(n9024), .B(n10431), .C(n7902), .Y(n3598) );
  OAI21X1 U1156 ( .A(n8983), .B(n10429), .C(n6287), .Y(n3599) );
  OAI21X1 U1158 ( .A(n9024), .B(n10428), .C(n6197), .Y(n3600) );
  OAI21X1 U1161 ( .A(n8983), .B(n10427), .C(n6196), .Y(n3601) );
  OAI21X1 U1163 ( .A(n9024), .B(n10426), .C(n7483), .Y(n3602) );
  OAI21X1 U1166 ( .A(n8983), .B(n10423), .C(n6121), .Y(n3603) );
  OAI21X1 U1168 ( .A(n9023), .B(n10422), .C(n7302), .Y(n3604) );
  OAI21X1 U1171 ( .A(n8983), .B(n10421), .C(n6056), .Y(n3605) );
  OAI21X1 U1173 ( .A(n9023), .B(n10420), .C(n7138), .Y(n3606) );
  OAI21X1 U1176 ( .A(n8982), .B(n10418), .C(n5112), .Y(n3607) );
  OAI21X1 U1178 ( .A(n9023), .B(n10417), .C(n6849), .Y(n3608) );
  OAI21X1 U1181 ( .A(n8982), .B(n10416), .C(n5111), .Y(n3609) );
  OAI21X1 U1183 ( .A(n9023), .B(n10415), .C(n6722), .Y(n3610) );
  OAI21X1 U1186 ( .A(n8982), .B(n10412), .C(n5110), .Y(n3611) );
  OAI21X1 U1188 ( .A(n9023), .B(n10411), .C(n6605), .Y(n3612) );
  OAI21X1 U1191 ( .A(n8982), .B(n10410), .C(n7900), .Y(n3613) );
  OAI21X1 U1193 ( .A(n9023), .B(n10409), .C(n6493), .Y(n3614) );
  OAI21X1 U1196 ( .A(n8982), .B(n10408), .C(n7685), .Y(n3615) );
  OAI21X1 U1198 ( .A(n9023), .B(n10407), .C(n7899), .Y(n3616) );
  OAI21X1 U1201 ( .A(n8982), .B(n10406), .C(n7481), .Y(n3617) );
  OAI21X1 U1203 ( .A(n9023), .B(n10405), .C(n8151), .Y(n3618) );
  OAI21X1 U1206 ( .A(n8982), .B(n10402), .C(n7301), .Y(n3619) );
  OAI21X1 U1208 ( .A(n9023), .B(n10401), .C(n7684), .Y(n3620) );
  OAI21X1 U1211 ( .A(n8982), .B(n10400), .C(n7137), .Y(n3621) );
  OAI21X1 U1213 ( .A(n9023), .B(n10399), .C(n7480), .Y(n3622) );
  OAI21X1 U1216 ( .A(n8982), .B(n10397), .C(n6989), .Y(n3623) );
  OAI21X1 U1218 ( .A(n9023), .B(n10396), .C(n6988), .Y(n3624) );
  OAI21X1 U1221 ( .A(n8981), .B(n10395), .C(n6848), .Y(n3625) );
  OAI21X1 U1223 ( .A(n9022), .B(n10394), .C(n7299), .Y(n3626) );
  OAI21X1 U1226 ( .A(n8981), .B(n10391), .C(n6604), .Y(n3627) );
  OAI21X1 U1228 ( .A(n9022), .B(n10390), .C(n7135), .Y(n3628) );
  OAI21X1 U1231 ( .A(n8981), .B(n10389), .C(n6492), .Y(n3629) );
  OAI21X1 U1233 ( .A(n9022), .B(n10388), .C(n6847), .Y(n3630) );
  OAI21X1 U1236 ( .A(n8987), .B(n10385), .C(n6721), .Y(n3631) );
  OAI21X1 U1238 ( .A(n9022), .B(n10384), .C(n6720), .Y(n3632) );
  OAI21X1 U1241 ( .A(n8981), .B(n10383), .C(n6386), .Y(n3633) );
  OAI21X1 U1243 ( .A(n9022), .B(n10382), .C(n6603), .Y(n3634) );
  OAI21X1 U1246 ( .A(n8982), .B(n10380), .C(n6285), .Y(n3635) );
  OAI21X1 U1248 ( .A(n9022), .B(n10379), .C(n6491), .Y(n3636) );
  OAI21X1 U1251 ( .A(n8982), .B(n10378), .C(n8149), .Y(n3637) );
  OAI21X1 U1253 ( .A(n9022), .B(n10377), .C(n8148), .Y(n3638) );
  OAI21X1 U1256 ( .A(n8982), .B(n10376), .C(n6845), .Y(n3639) );
  OAI21X1 U1258 ( .A(n9022), .B(n10375), .C(n6986), .Y(n3640) );
  OAI21X1 U1261 ( .A(n8982), .B(n10374), .C(n6718), .Y(n3641) );
  OAI21X1 U1263 ( .A(n9022), .B(n10373), .C(n6384), .Y(n3642) );
  OAI21X1 U1266 ( .A(n8982), .B(n10371), .C(n6601), .Y(n3643) );
  OAI21X1 U1268 ( .A(n9022), .B(n10370), .C(n6283), .Y(n3644) );
  OAI21X1 U1271 ( .A(n8983), .B(n10369), .C(n7898), .Y(n3645) );
  OAI21X1 U1273 ( .A(n8983), .B(n10366), .C(n7682), .Y(n3646) );
  OAI21X1 U1275 ( .A(n9022), .B(n10368), .C(n6193), .Y(n3647) );
  OAI21X1 U1278 ( .A(ap_CS_fsm[7]), .B(n10364), .C(n7897), .Y(n3648) );
  OAI21X1 U1281 ( .A(n9017), .B(n10363), .C(n8306), .Y(n3649) );
  OAI21X1 U1286 ( .A(n9012), .B(n10362), .C(n7681), .Y(n3651) );
  OAI21X1 U1289 ( .A(n9016), .B(n10361), .C(n8062), .Y(n3652) );
  OAI21X1 U1294 ( .A(ap_CS_fsm[7]), .B(n10360), .C(n7478), .Y(n3654) );
  OAI21X1 U1297 ( .A(n9015), .B(n10359), .C(n7840), .Y(n3655) );
  OAI21X1 U1302 ( .A(n9012), .B(n10358), .C(n7298), .Y(n3657) );
  OAI21X1 U1305 ( .A(n9016), .B(n10357), .C(n7628), .Y(n3658) );
  OAI21X1 U1311 ( .A(n6682), .B(n6683), .C(n9019), .Y(n1230) );
  NAND3X1 U1312 ( .A(n10270), .B(n1234), .C(n1235), .Y(n1232) );
  NOR3X1 U1313 ( .A(n7427), .B(n7425), .C(n7426), .Y(n1235) );
  NAND3X1 U1316 ( .A(n10257), .B(n10256), .C(n8257), .Y(n1236) );
  NOR3X1 U1318 ( .A(n7088), .B(CircularBuffer_head_i_read_ass_1_fu_1110_p3[10]), .C(n10271), .Y(n1234) );
  NAND3X1 U1321 ( .A(n1250), .B(tmp_33_i1_fu_1099_p2[3]), .C(
        tmp_33_i1_fu_1099_p2[4]), .Y(n1249) );
  NAND3X1 U1323 ( .A(n1251), .B(n1252), .C(n1253), .Y(n1231) );
  NOR3X1 U1324 ( .A(n7251), .B(n7249), .C(n7250), .Y(n1253) );
  NAND3X1 U1327 ( .A(n10268), .B(n10267), .C(n8256), .Y(n1254) );
  NOR3X1 U1329 ( .A(n6937), .B(CircularBuffer_head_i_read_ass_1_fu_1110_p3[26]), .C(CircularBuffer_head_i_read_ass_1_fu_1110_p3[25]), .Y(n1252) );
  NOR3X1 U1331 ( .A(n6806), .B(CircularBuffer_head_i_read_ass_1_fu_1110_p3[22]), .C(CircularBuffer_head_i_read_ass_1_fu_1110_p3[21]), .Y(n1251) );
  OAI21X1 U1333 ( .A(n9022), .B(n8661), .C(n6119), .Y(n3660) );
  OAI21X1 U1335 ( .A(n9020), .B(n8661), .C(n6844), .Y(n3661) );
  OAI21X1 U1338 ( .A(n9020), .B(n10244), .C(n6717), .Y(n3662) );
  OAI21X1 U1340 ( .A(n9020), .B(n10244), .C(n6600), .Y(n3663) );
  OAI21X1 U1343 ( .A(n9020), .B(n10245), .C(n8147), .Y(n3664) );
  OAI21X1 U1345 ( .A(n9020), .B(n10245), .C(n7477), .Y(n3665) );
  OAI21X1 U1348 ( .A(n9020), .B(n10246), .C(n7896), .Y(n3666) );
  OAI21X1 U1350 ( .A(n9020), .B(n10246), .C(n7297), .Y(n3667) );
  OAI21X1 U1353 ( .A(n9020), .B(n10247), .C(n7134), .Y(n3668) );
  OAI21X1 U1355 ( .A(n9020), .B(n10247), .C(n6985), .Y(n3669) );
  OAI21X1 U1358 ( .A(n9027), .B(n10248), .C(n6843), .Y(n3670) );
  OAI21X1 U1360 ( .A(n9023), .B(n10248), .C(n6489), .Y(n3671) );
  OAI21X1 U1363 ( .A(n9026), .B(n10249), .C(n6383), .Y(n3672) );
  OAI21X1 U1365 ( .A(n9029), .B(n10249), .C(n7680), .Y(n3673) );
  OAI21X1 U1368 ( .A(n9024), .B(n10250), .C(n6599), .Y(n3674) );
  OAI21X1 U1370 ( .A(n9025), .B(n10250), .C(n8146), .Y(n3675) );
  OAI21X1 U1373 ( .A(n9021), .B(n10251), .C(n7895), .Y(n3676) );
  OAI21X1 U1375 ( .A(n9022), .B(n10251), .C(n7476), .Y(n3677) );
  OAI21X1 U1378 ( .A(n9027), .B(n10252), .C(n7296), .Y(n3678) );
  OAI21X1 U1380 ( .A(n9028), .B(n10252), .C(n7133), .Y(n3679) );
  OAI21X1 U1383 ( .A(n9030), .B(n10253), .C(n6984), .Y(n3680) );
  OAI21X1 U1385 ( .A(n9020), .B(n10253), .C(n6842), .Y(n3681) );
  OAI21X1 U1388 ( .A(n9040), .B(n10254), .C(n6716), .Y(n3682) );
  OAI21X1 U1390 ( .A(n9023), .B(n10254), .C(n6488), .Y(n3683) );
  OAI21X1 U1393 ( .A(n9026), .B(n10255), .C(n6382), .Y(n3684) );
  OAI21X1 U1395 ( .A(n9021), .B(n10255), .C(n7679), .Y(n3685) );
  OAI21X1 U1398 ( .A(n9021), .B(n10256), .C(n6598), .Y(n3686) );
  OAI21X1 U1400 ( .A(n9021), .B(n10256), .C(n7894), .Y(n3687) );
  OAI21X1 U1403 ( .A(n9021), .B(n10257), .C(n7475), .Y(n3688) );
  OAI21X1 U1405 ( .A(n9021), .B(n10257), .C(n7132), .Y(n3689) );
  OAI21X1 U1408 ( .A(n9021), .B(n10258), .C(n6983), .Y(n3690) );
  OAI21X1 U1410 ( .A(n9021), .B(n10258), .C(n6841), .Y(n3691) );
  OAI21X1 U1413 ( .A(n9021), .B(n10259), .C(n6715), .Y(n3692) );
  OAI21X1 U1415 ( .A(n9021), .B(n10259), .C(n6487), .Y(n3693) );
  OAI21X1 U1418 ( .A(n9021), .B(n10260), .C(n6381), .Y(n3694) );
  OAI21X1 U1420 ( .A(n9021), .B(n10260), .C(n6282), .Y(n3695) );
  OAI21X1 U1423 ( .A(n9023), .B(n10261), .C(n6281), .Y(n3696) );
  OAI21X1 U1425 ( .A(n9031), .B(n10261), .C(n8145), .Y(n3697) );
  OAI21X1 U1428 ( .A(n9031), .B(n10262), .C(n7678), .Y(n3698) );
  OAI21X1 U1430 ( .A(n9031), .B(n10262), .C(n6192), .Y(n3699) );
  OAI21X1 U1433 ( .A(n9030), .B(n10263), .C(n7295), .Y(n3700) );
  OAI21X1 U1435 ( .A(n9030), .B(n10263), .C(n6280), .Y(n3701) );
  OAI21X1 U1438 ( .A(n9031), .B(n10264), .C(n6118), .Y(n3702) );
  OAI21X1 U1440 ( .A(n9030), .B(n10264), .C(n6191), .Y(n3703) );
  OAI21X1 U1443 ( .A(n9030), .B(n10265), .C(n6054), .Y(n3704) );
  OAI21X1 U1445 ( .A(n9030), .B(n10265), .C(n5109), .Y(n3705) );
  OAI21X1 U1448 ( .A(n9030), .B(n10266), .C(n6714), .Y(n3706) );
  OAI21X1 U1450 ( .A(n9030), .B(n10266), .C(n6117), .Y(n3707) );
  OAI21X1 U1453 ( .A(n9029), .B(n10267), .C(n6279), .Y(n3708) );
  OAI21X1 U1455 ( .A(n9029), .B(n10267), .C(n6190), .Y(n3709) );
  OAI21X1 U1458 ( .A(n9029), .B(n10268), .C(n6053), .Y(n3710) );
  OAI21X1 U1460 ( .A(n9029), .B(n10268), .C(n5108), .Y(n3711) );
  OAI21X1 U1463 ( .A(n9029), .B(n10269), .C(n6486), .Y(n3712) );
  OAI21X1 U1465 ( .A(n9029), .B(n10269), .C(n5107), .Y(n3713) );
  OAI21X1 U1468 ( .A(n9028), .B(recentABools_head_i[0]), .C(n6052), .Y(n3714)
         );
  OAI21X1 U1471 ( .A(n9012), .B(n10272), .C(n6982), .Y(n3715) );
  OAI21X1 U1474 ( .A(n9016), .B(n10271), .C(n6189), .Y(n3716) );
  OAI21X1 U1477 ( .A(n9028), .B(n8662), .C(n7131), .Y(n3717) );
  OAI21X1 U1479 ( .A(n9028), .B(n8430), .C(n6380), .Y(n3718) );
  OAI21X1 U1481 ( .A(n9028), .B(n8431), .C(n6278), .Y(n3719) );
  OAI21X1 U1483 ( .A(n9028), .B(n8432), .C(n6188), .Y(n3720) );
  OAI21X1 U1485 ( .A(n9028), .B(n8433), .C(n6116), .Y(n3721) );
  OAI21X1 U1487 ( .A(n9028), .B(n8434), .C(n5106), .Y(n3722) );
  OAI21X1 U1489 ( .A(n9027), .B(n8435), .C(n6051), .Y(n3723) );
  OAI21X1 U1491 ( .A(n9027), .B(n8436), .C(n6379), .Y(n3724) );
  OAI21X1 U1493 ( .A(n9027), .B(n8437), .C(n6115), .Y(n3725) );
  OAI21X1 U1495 ( .A(n9030), .B(n8438), .C(n5105), .Y(n3726) );
  OAI21X1 U1497 ( .A(n9027), .B(n8439), .C(n5104), .Y(n3727) );
  OAI21X1 U1499 ( .A(n9027), .B(n8440), .C(n6981), .Y(n3728) );
  OAI21X1 U1501 ( .A(n9027), .B(n8441), .C(n6597), .Y(n3729) );
  OAI21X1 U1503 ( .A(n9028), .B(n8442), .C(n5103), .Y(n3730) );
  OAI21X1 U1505 ( .A(n9028), .B(n8443), .C(n5102), .Y(n3731) );
  OAI21X1 U1507 ( .A(n9028), .B(n8444), .C(n5101), .Y(n3732) );
  OAI21X1 U1509 ( .A(n9028), .B(n8445), .C(n5100), .Y(n3733) );
  OAI21X1 U1511 ( .A(n9028), .B(n8446), .C(n5099), .Y(n3734) );
  OAI21X1 U1513 ( .A(n9029), .B(n8447), .C(n6114), .Y(n3735) );
  OAI21X1 U1515 ( .A(n9029), .B(n8448), .C(n5098), .Y(n3736) );
  OAI21X1 U1517 ( .A(n9029), .B(n8449), .C(n6378), .Y(n3737) );
  OAI21X1 U1519 ( .A(n9029), .B(n8450), .C(n5097), .Y(n3738) );
  OAI21X1 U1521 ( .A(n9029), .B(n8451), .C(n5096), .Y(n3739) );
  OAI21X1 U1523 ( .A(n9029), .B(n8452), .C(n7893), .Y(n3740) );
  OAI21X1 U1525 ( .A(n9030), .B(n8453), .C(n7474), .Y(n3741) );
  OAI21X1 U1527 ( .A(n9030), .B(n8454), .C(n7130), .Y(n3742) );
  OAI21X1 U1529 ( .A(n9031), .B(n8455), .C(n6277), .Y(n3743) );
  OAI21X1 U1531 ( .A(n9030), .B(n8456), .C(n5095), .Y(n3744) );
  OAI21X1 U1533 ( .A(n9031), .B(n8457), .C(n6050), .Y(n3745) );
  OAI21X1 U1535 ( .A(n9030), .B(n8458), .C(n5094), .Y(n3746) );
  OAI21X1 U1537 ( .A(n9031), .B(n8489), .C(n5093), .Y(n3747) );
  AOI22X1 U1540 ( .A(N496), .B(ap_CS_fsm[8]), .C(\tmp_12_reg_1694[0] ), .D(
        n10242), .Y(n1401) );
  OAI21X1 U1542 ( .A(n9004), .B(n4688), .C(n7673), .Y(n3749) );
  OAI21X1 U1544 ( .A(n9005), .B(n8459), .C(n8141), .Y(n3750) );
  OAI21X1 U1546 ( .A(n9005), .B(n8460), .C(n7888), .Y(n3751) );
  OAI21X1 U1548 ( .A(n9005), .B(n8461), .C(n7672), .Y(n3752) );
  OAI21X1 U1550 ( .A(n9004), .B(n8462), .C(n7468), .Y(n3753) );
  OAI21X1 U1552 ( .A(n9004), .B(n8463), .C(n8140), .Y(n3754) );
  OAI21X1 U1554 ( .A(n9004), .B(n8464), .C(n7887), .Y(n3755) );
  OAI21X1 U1556 ( .A(n9004), .B(n8465), .C(n7289), .Y(n3756) );
  OAI21X1 U1558 ( .A(n9003), .B(n8466), .C(n7467), .Y(n3757) );
  OAI21X1 U1560 ( .A(n9003), .B(n8467), .C(n7288), .Y(n3758) );
  OAI21X1 U1562 ( .A(n9003), .B(n8468), .C(n7124), .Y(n3759) );
  OAI21X1 U1564 ( .A(n9002), .B(n8469), .C(n6975), .Y(n3760) );
  OAI21X1 U1566 ( .A(n9002), .B(n8470), .C(n7466), .Y(n3761) );
  OAI21X1 U1568 ( .A(n9002), .B(n8471), .C(n7287), .Y(n3762) );
  OAI21X1 U1570 ( .A(n9002), .B(n8472), .C(n6836), .Y(n3763) );
  OAI21X1 U1572 ( .A(n9001), .B(n8473), .C(n6974), .Y(n3764) );
  OAI21X1 U1574 ( .A(n9001), .B(n8474), .C(n6709), .Y(n3765) );
  OAI21X1 U1576 ( .A(n9001), .B(n8475), .C(n6592), .Y(n3766) );
  OAI21X1 U1578 ( .A(n9001), .B(n8476), .C(n6481), .Y(n3767) );
  OAI21X1 U1580 ( .A(n9000), .B(n8477), .C(n7123), .Y(n3768) );
  OAI21X1 U1582 ( .A(n9000), .B(n8478), .C(n6835), .Y(n3769) );
  OAI21X1 U1584 ( .A(n9000), .B(n8479), .C(n6373), .Y(n3770) );
  OAI21X1 U1586 ( .A(n9000), .B(n8480), .C(n6272), .Y(n3771) );
  OAI21X1 U1588 ( .A(n8999), .B(n8481), .C(n6183), .Y(n3772) );
  OAI21X1 U1590 ( .A(n8999), .B(n8482), .C(n6109), .Y(n3773) );
  OAI21X1 U1592 ( .A(n8999), .B(n8483), .C(n6708), .Y(n3774) );
  OAI21X1 U1594 ( .A(n8999), .B(n8484), .C(n6591), .Y(n3775) );
  OAI21X1 U1596 ( .A(n8998), .B(n8485), .C(n6480), .Y(n3776) );
  OAI21X1 U1598 ( .A(n8998), .B(n8486), .C(n6372), .Y(n3777) );
  OAI21X1 U1600 ( .A(n8998), .B(n8487), .C(n6271), .Y(n3778) );
  OAI21X1 U1602 ( .A(n8998), .B(n8488), .C(n6182), .Y(n3779) );
  OAI21X1 U1604 ( .A(n9002), .B(n8663), .C(n8139), .Y(n3780) );
  OAI21X1 U1606 ( .A(n11046), .B(n1468), .C(n7077), .Y(n3781) );
  OAI21X1 U1608 ( .A(n7078), .B(n7233), .C(ap_CS_fsm[6]), .Y(n1468) );
  NAND3X1 U1609 ( .A(n1473), .B(n1474), .C(n1475), .Y(n1472) );
  NOR3X1 U1610 ( .A(n8274), .B(n7802), .C(n8038), .Y(n1475) );
  NAND3X1 U1613 ( .A(n10098), .B(n10099), .C(n8275), .Y(n1476) );
  NOR3X1 U1615 ( .A(n7600), .B(CircularBuffer_len_read_assign_1_reg_1616[14]), 
        .C(CircularBuffer_len_read_assign_1_reg_1616[13]), .Y(n1474) );
  NOR3X1 U1617 ( .A(n7409), .B(CircularBuffer_len_read_assign_1_reg_1616[10]), 
        .C(CircularBuffer_len_write_assig_1_fu_924_p2[0]), .Y(n1473) );
  NAND3X1 U1619 ( .A(n1492), .B(n1493), .C(n1494), .Y(n1471) );
  NOR3X1 U1620 ( .A(n8025), .B(n8023), .C(n8024), .Y(n1494) );
  NAND3X1 U1623 ( .A(n10084), .B(n10085), .C(n8251), .Y(n1495) );
  NOR3X1 U1625 ( .A(n7799), .B(CircularBuffer_len_read_assign_1_reg_1616[29]), 
        .C(CircularBuffer_len_read_assign_1_reg_1616[28]), .Y(n1493) );
  NOR3X1 U1627 ( .A(n8270), .B(CircularBuffer_len_read_assign_1_reg_1616[25]), 
        .C(CircularBuffer_len_read_assign_1_reg_1616[24]), .Y(n1492) );
  OAI21X1 U1629 ( .A(n11046), .B(n9934), .C(n8138), .Y(n3782) );
  NAND3X1 U1633 ( .A(\not_tmp_i_i4_reg_1650[0] ), .B(ap_CS_fsm[6]), .C(
        \recentVBools_data_q1[0] ), .Y(n1514) );
  AOI22X1 U1636 ( .A(N513), .B(ap_CS_fsm[3]), .C(\tmp_s_reg_1578[0] ), .D(
        n9934), .Y(n1515) );
  AOI22X1 U1638 ( .A(n1516), .B(n1517), .C(n10056), .D(n10171), .Y(n3785) );
  NOR3X1 U1640 ( .A(n7235), .B(n7606), .C(n8043), .Y(n1517) );
  NAND3X1 U1641 ( .A(n10162), .B(n10163), .C(n8044), .Y(n1522) );
  NAND3X1 U1643 ( .A(n10166), .B(n10167), .C(n7607), .Y(n1521) );
  NOR3X1 U1646 ( .A(n7236), .B(CircularBuffer_len_write_assig_reg_1634[6]), 
        .C(CircularBuffer_len_write_assig_reg_1634[5]), .Y(n1530) );
  NAND3X1 U1647 ( .A(n10147), .B(n10148), .C(n10146), .Y(n1531) );
  NOR3X1 U1648 ( .A(n8280), .B(CircularBuffer_len_write_assig_reg_1634[31]), 
        .C(CircularBuffer_len_write_assig_reg_1634[30]), .Y(n1529) );
  NOR3X1 U1650 ( .A(n7411), .B(n7806), .C(n8286), .Y(n1516) );
  NAND3X1 U1651 ( .A(n10155), .B(n10156), .C(n8287), .Y(n1540) );
  NAND3X1 U1653 ( .A(n10140), .B(n10159), .C(n7807), .Y(n1539) );
  NOR3X1 U1656 ( .A(n7412), .B(CircularBuffer_len_write_assig_reg_1634[13]), 
        .C(CircularBuffer_len_write_assig_reg_1634[12]), .Y(n1548) );
  NOR3X1 U1658 ( .A(n8272), .B(CircularBuffer_len_write_assig_reg_1634[11]), 
        .C(CircularBuffer_len_write_assig_reg_1634[10]), .Y(n1547) );
  OAI21X1 U1660 ( .A(n8894), .B(n10170), .C(n5092), .Y(n3786) );
  OAI21X1 U1663 ( .A(n8894), .B(n10169), .C(n7886), .Y(n3787) );
  OAI21X1 U1666 ( .A(n8894), .B(n10168), .C(n5091), .Y(n3788) );
  OAI21X1 U1669 ( .A(n1646), .B(n10167), .C(n5090), .Y(n3789) );
  OAI21X1 U1672 ( .A(n8894), .B(n10166), .C(n5089), .Y(n3790) );
  OAI21X1 U1675 ( .A(n1646), .B(n10165), .C(n5088), .Y(n3791) );
  OAI21X1 U1678 ( .A(n1646), .B(n10164), .C(n5087), .Y(n3792) );
  OAI21X1 U1681 ( .A(n8894), .B(n10163), .C(n5086), .Y(n3793) );
  OAI21X1 U1684 ( .A(n1646), .B(n10162), .C(n7465), .Y(n3794) );
  OAI21X1 U1687 ( .A(n8894), .B(n10161), .C(n5085), .Y(n3795) );
  OAI21X1 U1690 ( .A(n1646), .B(n10160), .C(n5084), .Y(n3796) );
  OAI21X1 U1693 ( .A(n1646), .B(n10159), .C(n5083), .Y(n3797) );
  OAI21X1 U1696 ( .A(n1646), .B(n10158), .C(n5082), .Y(n3798) );
  OAI21X1 U1699 ( .A(n8894), .B(n10157), .C(n5081), .Y(n3799) );
  OAI21X1 U1702 ( .A(n1646), .B(n10156), .C(n5080), .Y(n3800) );
  OAI21X1 U1705 ( .A(n8894), .B(n10155), .C(n5079), .Y(n3801) );
  OAI21X1 U1708 ( .A(n8894), .B(n10154), .C(n6973), .Y(n3802) );
  OAI21X1 U1711 ( .A(n1646), .B(n10153), .C(n6834), .Y(n3803) );
  OAI21X1 U1714 ( .A(n1646), .B(n10152), .C(n5078), .Y(n3804) );
  OAI21X1 U1717 ( .A(n8894), .B(n10151), .C(n5077), .Y(n3805) );
  OAI21X1 U1720 ( .A(n1646), .B(n10150), .C(n7558), .Y(n3806) );
  OAI21X1 U1723 ( .A(n1646), .B(n10149), .C(n7217), .Y(n3807) );
  OAI21X1 U1726 ( .A(n1646), .B(n10148), .C(n7286), .Y(n3808) );
  OAI21X1 U1729 ( .A(n1646), .B(n10147), .C(n7669), .Y(n3809) );
  OAI21X1 U1732 ( .A(n8894), .B(n10146), .C(n6707), .Y(n3810) );
  OAI21X1 U1735 ( .A(n1646), .B(n10145), .C(n5076), .Y(n3811) );
  OAI21X1 U1738 ( .A(n1646), .B(n10144), .C(n6972), .Y(n3812) );
  OAI21X1 U1741 ( .A(n1646), .B(n10143), .C(n6833), .Y(n3813) );
  OAI21X1 U1744 ( .A(n8894), .B(n10142), .C(n6706), .Y(n3814) );
  OAI21X1 U1747 ( .A(n8894), .B(n10141), .C(n6590), .Y(n3815) );
  OAI21X1 U1750 ( .A(n1646), .B(n10140), .C(n6479), .Y(n3816) );
  OAI21X1 U1753 ( .A(n1646), .B(n10139), .C(n6371), .Y(n3817) );
  OAI21X1 U1756 ( .A(n8983), .B(n10109), .C(n7461), .Y(n3818) );
  OAI21X1 U1759 ( .A(n8983), .B(n10108), .C(n8134), .Y(n3819) );
  OAI21X1 U1762 ( .A(n8983), .B(n10107), .C(n5075), .Y(n3820) );
  OAI21X1 U1765 ( .A(n8984), .B(n10106), .C(n5074), .Y(n3821) );
  OAI21X1 U1768 ( .A(n8984), .B(n10105), .C(n6700), .Y(n3822) );
  OAI21X1 U1771 ( .A(n8984), .B(n10104), .C(n6585), .Y(n3823) );
  OAI21X1 U1774 ( .A(n8984), .B(n10103), .C(n6366), .Y(n3824) );
  OAI21X1 U1777 ( .A(n8985), .B(n10102), .C(n5073), .Y(n3825) );
  OAI21X1 U1780 ( .A(n8985), .B(n10101), .C(n7282), .Y(n3826) );
  OAI21X1 U1783 ( .A(n8985), .B(n10100), .C(n5072), .Y(n3827) );
  OAI21X1 U1786 ( .A(n8985), .B(n10099), .C(n5071), .Y(n3828) );
  OAI21X1 U1789 ( .A(n8985), .B(n10098), .C(n5070), .Y(n3829) );
  OAI21X1 U1792 ( .A(n8986), .B(n10097), .C(n6474), .Y(n3830) );
  OAI21X1 U1795 ( .A(n8986), .B(n10096), .C(n6365), .Y(n3831) );
  OAI21X1 U1798 ( .A(n8986), .B(n10095), .C(n6179), .Y(n3832) );
  OAI21X1 U1801 ( .A(n8986), .B(n10094), .C(n6106), .Y(n3833) );
  OAI21X1 U1804 ( .A(n8986), .B(n10093), .C(n6046), .Y(n3834) );
  OAI21X1 U1807 ( .A(n8991), .B(n10092), .C(n6967), .Y(n3835) );
  OAI21X1 U1810 ( .A(n8990), .B(n10091), .C(n7281), .Y(n3836) );
  OAI21X1 U1813 ( .A(n8990), .B(n10090), .C(n7118), .Y(n3837) );
  OAI21X1 U1816 ( .A(n8990), .B(n10089), .C(n6045), .Y(n3838) );
  OAI21X1 U1819 ( .A(n8990), .B(n10088), .C(n6828), .Y(n3839) );
  OAI21X1 U1822 ( .A(n8990), .B(n10087), .C(n5069), .Y(n3840) );
  OAI21X1 U1825 ( .A(n8989), .B(n10086), .C(n6266), .Y(n3841) );
  OAI21X1 U1828 ( .A(n8989), .B(n10085), .C(n6178), .Y(n3842) );
  OAI21X1 U1831 ( .A(n8989), .B(n10084), .C(n6105), .Y(n3843) );
  OAI21X1 U1834 ( .A(n8989), .B(n10083), .C(n5068), .Y(n3844) );
  OAI21X1 U1837 ( .A(n8988), .B(n10082), .C(n7117), .Y(n3845) );
  OAI21X1 U1840 ( .A(n8988), .B(n10081), .C(n5067), .Y(n3846) );
  OAI21X1 U1843 ( .A(n8988), .B(n10080), .C(n7883), .Y(n3847) );
  OAI21X1 U1846 ( .A(n8988), .B(n10079), .C(n5066), .Y(n3848) );
  OAI21X1 U1849 ( .A(n8987), .B(n10077), .C(n8895), .Y(n3849) );
  OAI21X1 U1851 ( .A(n8987), .B(n10076), .C(n6104), .Y(n3850) );
  OAI21X1 U1854 ( .A(n5548), .B(n5718), .C(n5065), .Y(n3851) );
  NAND3X1 U1856 ( .A(n1652), .B(n1653), .C(n1654), .Y(n1650) );
  NOR3X1 U1857 ( .A(n8042), .B(n8040), .C(n8041), .Y(n1654) );
  NAND3X1 U1860 ( .A(n9914), .B(n9913), .C(n8250), .Y(n1655) );
  NOR3X1 U1862 ( .A(n8269), .B(tmp_38_i_reg_1550[11]), .C(
        tmp_38_i_reg_1550[10]), .Y(n1653) );
  NOR3X1 U1864 ( .A(n7798), .B(n9830), .C(n9928), .Y(n1652) );
  NAND3X1 U1866 ( .A(n1672), .B(n1673), .C(n1674), .Y(n1649) );
  NOR3X1 U1867 ( .A(n5895), .B(n5899), .C(n5905), .Y(n1674) );
  NAND3X1 U1869 ( .A(n9924), .B(n9923), .C(n9925), .Y(n1676) );
  NAND3X1 U1870 ( .A(n9903), .B(n9902), .C(n8264), .Y(n1675) );
  NOR3X1 U1872 ( .A(n7408), .B(tmp_38_i_reg_1550[26]), .C(
        tmp_38_i_reg_1550[25]), .Y(n1673) );
  NOR3X1 U1874 ( .A(n7599), .B(tmp_38_i_reg_1550[22]), .C(
        tmp_38_i_reg_1550[21]), .Y(n1672) );
  OAI21X1 U1876 ( .A(ap_CS_fsm[2]), .B(n10055), .C(n8133), .Y(n3852) );
  OAI21X1 U1879 ( .A(n8987), .B(n10054), .C(n8305), .Y(n3853) );
  OAI21X1 U1884 ( .A(ap_CS_fsm[2]), .B(n10053), .C(n7882), .Y(n3855) );
  OAI21X1 U1887 ( .A(n8987), .B(n10052), .C(n8061), .Y(n3856) );
  OAI21X1 U1894 ( .A(ap_CS_fsm[2]), .B(n10051), .C(n7667), .Y(n3859) );
  OAI21X1 U1897 ( .A(n8987), .B(n10050), .C(n7839), .Y(n3860) );
  OAI21X1 U1902 ( .A(n8998), .B(n8660), .C(n6966), .Y(n3862) );
  OAI21X1 U1904 ( .A(n8998), .B(n8660), .C(n6827), .Y(n3863) );
  OAI21X1 U1906 ( .A(n8999), .B(n9936), .C(n6473), .Y(n3864) );
  OAI21X1 U1908 ( .A(n8999), .B(n9936), .C(n6363), .Y(n3865) );
  OAI21X1 U1910 ( .A(n8999), .B(n9937), .C(n6265), .Y(n3866) );
  OAI21X1 U1912 ( .A(n8999), .B(n9937), .C(n6044), .Y(n3867) );
  OAI21X1 U1914 ( .A(n8999), .B(n9938), .C(n7116), .Y(n3868) );
  OAI21X1 U1916 ( .A(n8999), .B(n9938), .C(n5064), .Y(n3869) );
  OAI21X1 U1918 ( .A(n8999), .B(n9939), .C(n5063), .Y(n3870) );
  OAI21X1 U1920 ( .A(n8999), .B(n9939), .C(n5062), .Y(n3871) );
  OAI21X1 U1922 ( .A(n9000), .B(n9940), .C(n8132), .Y(n3872) );
  OAI21X1 U1924 ( .A(n9000), .B(n9940), .C(n7666), .Y(n3873) );
  OAI21X1 U1927 ( .A(n9000), .B(n9941), .C(n7881), .Y(n3874) );
  OAI21X1 U1929 ( .A(n9000), .B(n9941), .C(n7460), .Y(n3875) );
  OAI21X1 U1932 ( .A(n9000), .B(n9942), .C(n7280), .Y(n3876) );
  OAI21X1 U1934 ( .A(n9000), .B(n9942), .C(n6965), .Y(n3877) );
  OAI21X1 U1936 ( .A(n9000), .B(n9943), .C(n6584), .Y(n3878) );
  OAI21X1 U1938 ( .A(n9000), .B(n9943), .C(n6472), .Y(n3879) );
  OAI21X1 U1940 ( .A(n9001), .B(n9944), .C(n7115), .Y(n3880) );
  OAI21X1 U1942 ( .A(n9001), .B(n9944), .C(n6826), .Y(n3881) );
  OAI21X1 U1945 ( .A(n9001), .B(n9945), .C(n6362), .Y(n3882) );
  OAI21X1 U1947 ( .A(n9001), .B(n9945), .C(n6264), .Y(n3883) );
  OAI21X1 U1950 ( .A(n9001), .B(n9946), .C(n6176), .Y(n3884) );
  OAI21X1 U1952 ( .A(n9001), .B(n9946), .C(n6103), .Y(n3885) );
  OAI21X1 U1955 ( .A(n9001), .B(n9947), .C(n6043), .Y(n3886) );
  OAI21X1 U1957 ( .A(n9001), .B(n9947), .C(n8131), .Y(n3887) );
  OAI21X1 U1960 ( .A(n9002), .B(n9948), .C(n7880), .Y(n3888) );
  OAI21X1 U1962 ( .A(n9002), .B(n9948), .C(n7665), .Y(n3889) );
  OAI21X1 U1964 ( .A(n9002), .B(n9949), .C(n7114), .Y(n3890) );
  OAI21X1 U1966 ( .A(n9002), .B(n9949), .C(n6699), .Y(n3891) );
  OAI21X1 U1968 ( .A(n9002), .B(n9950), .C(n6583), .Y(n3892) );
  OAI21X1 U1970 ( .A(n9002), .B(n9950), .C(n6471), .Y(n3893) );
  OAI21X1 U1972 ( .A(n9002), .B(n9951), .C(n6361), .Y(n3894) );
  OAI21X1 U1974 ( .A(n9003), .B(n9951), .C(n6964), .Y(n3895) );
  OAI21X1 U1976 ( .A(n9003), .B(n9952), .C(n6825), .Y(n3896) );
  OAI21X1 U1978 ( .A(n9003), .B(n9952), .C(n6263), .Y(n3897) );
  OAI21X1 U1980 ( .A(n9003), .B(n9953), .C(n6175), .Y(n3898) );
  OAI21X1 U1982 ( .A(n9003), .B(n9953), .C(n6102), .Y(n3899) );
  OAI21X1 U1984 ( .A(n9003), .B(n9954), .C(n6042), .Y(n3900) );
  OAI21X1 U1986 ( .A(n9003), .B(n9954), .C(n5061), .Y(n3901) );
  OAI21X1 U1988 ( .A(n9003), .B(n9955), .C(n5060), .Y(n3902) );
  OAI21X1 U1990 ( .A(n9004), .B(n9955), .C(n7113), .Y(n3903) );
  OAI21X1 U1992 ( .A(n9004), .B(n9956), .C(n6963), .Y(n3904) );
  OAI21X1 U1994 ( .A(n9004), .B(n9956), .C(n6824), .Y(n3905) );
  OAI21X1 U1997 ( .A(n9004), .B(n9957), .C(n6698), .Y(n3906) );
  OAI21X1 U1999 ( .A(n9005), .B(n9957), .C(n6582), .Y(n3907) );
  OAI21X1 U2002 ( .A(n9003), .B(n9958), .C(n8130), .Y(n3908) );
  OAI21X1 U2004 ( .A(n9004), .B(n9958), .C(n6470), .Y(n3909) );
  OAI21X1 U2007 ( .A(n9005), .B(n9959), .C(n6360), .Y(n3910) );
  OAI21X1 U2009 ( .A(n9005), .B(n9959), .C(n6262), .Y(n3911) );
  OAI21X1 U2011 ( .A(n9005), .B(n9960), .C(n6174), .Y(n3912) );
  OAI21X1 U2013 ( .A(n9004), .B(n9960), .C(n6101), .Y(n3913) );
  OAI21X1 U2015 ( .A(n9005), .B(n9961), .C(n6041), .Y(n3914) );
  OAI21X1 U2017 ( .A(n9005), .B(n9961), .C(n5059), .Y(n3915) );
  OAI21X1 U2019 ( .A(ap_CS_fsm[2]), .B(n10025), .C(n7459), .Y(n3916) );
  OAI21X1 U2022 ( .A(n8987), .B(n10024), .C(n5058), .Y(n3917) );
  OAI21X1 U2025 ( .A(n9004), .B(recentVBools_head_i[0]), .C(n5057), .Y(n3918)
         );
  OAI21X1 U2028 ( .A(ap_CS_fsm[2]), .B(n9964), .C(n7279), .Y(n3919) );
  OAI21X1 U2031 ( .A(n8981), .B(n9963), .C(n7627), .Y(n3920) );
  OAI21X1 U2034 ( .A(n6680), .B(n6681), .C(ap_CS_fsm[4]), .Y(n1800) );
  NAND3X1 U2035 ( .A(n9962), .B(n1804), .C(n1805), .Y(n1802) );
  NOR3X1 U2036 ( .A(n7424), .B(n7422), .C(n7423), .Y(n1805) );
  NAND3X1 U2043 ( .A(n9949), .B(n9948), .C(n8255), .Y(n1806) );
  NOR3X1 U2047 ( .A(n7087), .B(CircularBuffer_head_i_read_ass_fu_797_p3[10]), 
        .C(n10024), .Y(n1804) );
  NAND3X1 U2052 ( .A(n1812), .B(tmp_33_i_fu_786_p2[3]), .C(
        tmp_33_i_fu_786_p2[4]), .Y(n1811) );
  NAND3X1 U2054 ( .A(n1813), .B(n1814), .C(n1815), .Y(n1801) );
  NOR3X1 U2055 ( .A(n7248), .B(n7246), .C(n7247), .Y(n1815) );
  NAND3X1 U2062 ( .A(n9960), .B(n9959), .C(n8254), .Y(n1816) );
  NOR3X1 U2066 ( .A(n6936), .B(CircularBuffer_head_i_read_ass_fu_797_p3[26]), 
        .C(CircularBuffer_head_i_read_ass_fu_797_p3[25]), .Y(n1814) );
  NOR3X1 U2070 ( .A(n6805), .B(CircularBuffer_head_i_read_ass_fu_797_p3[22]), 
        .C(CircularBuffer_head_i_read_ass_fu_797_p3[21]), .Y(n1813) );
  OAI21X1 U2075 ( .A(ap_CS_fsm[1]), .B(n9929), .C(n6684), .Y(n3921) );
  OAI21X1 U2076 ( .A(n8976), .B(n9928), .C(n8060), .Y(n3922) );
  OAI21X1 U2077 ( .A(n8975), .B(n9927), .C(n6808), .Y(n3923) );
  OAI21X1 U2078 ( .A(ap_CS_fsm[1]), .B(n9926), .C(n6941), .Y(n3924) );
  OAI21X1 U2079 ( .A(n8976), .B(n9925), .C(n7091), .Y(n3925) );
  OAI21X1 U2080 ( .A(n8975), .B(n9924), .C(n7255), .Y(n3926) );
  OAI21X1 U2082 ( .A(ap_CS_fsm[1]), .B(n9923), .C(n7431), .Y(n3927) );
  OAI21X1 U2084 ( .A(n8976), .B(n9922), .C(n6456), .Y(n3928) );
  OAI21X1 U2086 ( .A(n8975), .B(n9921), .C(n7622), .Y(n3929) );
  OAI21X1 U2087 ( .A(ap_CS_fsm[1]), .B(n9920), .C(n7835), .Y(n3930) );
  OAI21X1 U2088 ( .A(n8976), .B(n9919), .C(n8057), .Y(n3931) );
  OAI21X1 U2090 ( .A(n8975), .B(n9918), .C(n8300), .Y(n3932) );
  OAI21X1 U2092 ( .A(n8975), .B(n9917), .C(n6348), .Y(n3933) );
  OAI21X1 U2093 ( .A(n8976), .B(n9916), .C(n6457), .Y(n3934) );
  OAI21X1 U2094 ( .A(ap_CS_fsm[1]), .B(n9915), .C(n6570), .Y(n3935) );
  OAI21X1 U2095 ( .A(ap_CS_fsm[1]), .B(n9914), .C(n6685), .Y(n3936) );
  OAI21X1 U2096 ( .A(ap_CS_fsm[1]), .B(n9913), .C(n6809), .Y(n3937) );
  OAI21X1 U2097 ( .A(n8976), .B(n9912), .C(n6942), .Y(n3938) );
  OAI21X1 U2098 ( .A(n8975), .B(n9911), .C(n7092), .Y(n3939) );
  OAI21X1 U2099 ( .A(n8976), .B(n9910), .C(n7256), .Y(n3940) );
  OAI21X1 U2101 ( .A(n8976), .B(n9909), .C(n7432), .Y(n3941) );
  OAI21X1 U2103 ( .A(ap_CS_fsm[1]), .B(n9908), .C(n7623), .Y(n3942) );
  OAI21X1 U2105 ( .A(ap_CS_fsm[1]), .B(n9907), .C(n7836), .Y(n3943) );
  OAI21X1 U2107 ( .A(ap_CS_fsm[1]), .B(n9906), .C(n8058), .Y(n3944) );
  OAI21X1 U2108 ( .A(n8975), .B(n9905), .C(n8301), .Y(n3945) );
  OAI21X1 U2109 ( .A(n8975), .B(n9904), .C(n7624), .Y(n3946) );
  OAI21X1 U2111 ( .A(n8975), .B(n9903), .C(n7837), .Y(n3947) );
  OAI21X1 U2113 ( .A(n8975), .B(n9902), .C(n8059), .Y(n3948) );
  OAI21X1 U2114 ( .A(n8975), .B(n9901), .C(n8302), .Y(n3949) );
  OAI21X1 U2115 ( .A(n8975), .B(n9900), .C(n6943), .Y(n3950) );
  OAI21X1 U2117 ( .A(n8975), .B(n9899), .C(n7093), .Y(n3951) );
  OAI21X1 U2119 ( .A(n8975), .B(n9898), .C(n7626), .Y(n3952) );
  OAI21X1 U2121 ( .A(n8975), .B(n9897), .C(n7257), .Y(n3953) );
  OAI21X1 U2123 ( .A(n8975), .B(n9896), .C(n7433), .Y(n3954) );
  OAI21X1 U2125 ( .A(n8977), .B(n9885), .C(n8129), .Y(n3955) );
  OAI21X1 U2127 ( .A(n8977), .B(n9884), .C(n7879), .Y(n3956) );
  OAI21X1 U2129 ( .A(n8977), .B(n9883), .C(n7664), .Y(n3957) );
  OAI21X1 U2131 ( .A(n8977), .B(n9882), .C(n7458), .Y(n3958) );
  OAI21X1 U2133 ( .A(n8977), .B(n9881), .C(n7278), .Y(n3959) );
  OAI21X1 U2135 ( .A(n8977), .B(n9880), .C(n7112), .Y(n3960) );
  OAI21X1 U2137 ( .A(n8977), .B(n9879), .C(n6962), .Y(n3961) );
  OAI21X1 U2139 ( .A(n8977), .B(n9878), .C(n8128), .Y(n3962) );
  OAI21X1 U2141 ( .A(n8977), .B(n9877), .C(n6823), .Y(n3963) );
  OAI21X1 U2143 ( .A(n8977), .B(n9876), .C(n6697), .Y(n3964) );
  OAI21X1 U2145 ( .A(n8977), .B(n9875), .C(n6581), .Y(n3965) );
  OAI21X1 U2147 ( .A(n8977), .B(n9874), .C(n6469), .Y(n3966) );
  OAI21X1 U2149 ( .A(n8977), .B(n9873), .C(n6359), .Y(n3967) );
  OAI21X1 U2151 ( .A(n8977), .B(n9872), .C(n7878), .Y(n3968) );
  OAI21X1 U2153 ( .A(n8980), .B(n9871), .C(n7663), .Y(n3969) );
  OAI21X1 U2155 ( .A(n8979), .B(n9870), .C(n7277), .Y(n3970) );
  OAI21X1 U2157 ( .A(n8978), .B(n9869), .C(n6696), .Y(n3971) );
  OAI21X1 U2159 ( .A(n8977), .B(n9868), .C(n7457), .Y(n3972) );
  OAI21X1 U2161 ( .A(n8980), .B(n9867), .C(n7111), .Y(n3973) );
  OAI21X1 U2163 ( .A(n8979), .B(n9866), .C(n6961), .Y(n3974) );
  OAI21X1 U2165 ( .A(n8978), .B(n9865), .C(n6822), .Y(n3975) );
  OAI21X1 U2167 ( .A(n8978), .B(n9864), .C(n8127), .Y(n3976) );
  OAI21X1 U2169 ( .A(n8980), .B(n9863), .C(n6580), .Y(n3977) );
  OAI21X1 U2171 ( .A(n8979), .B(n9862), .C(n6468), .Y(n3978) );
  OAI21X1 U2173 ( .A(n8978), .B(n9861), .C(n6358), .Y(n3979) );
  OAI21X1 U2175 ( .A(n8980), .B(n9860), .C(n7877), .Y(n3980) );
  OAI21X1 U2177 ( .A(n8977), .B(n8659), .C(n6695), .Y(n3981) );
  OAI21X1 U2179 ( .A(n8962), .B(n9895), .C(n6467), .Y(n3982) );
  OAI21X1 U2182 ( .A(n8975), .B(n9894), .C(n7626), .Y(n3983) );
  NAND3X1 U2183 ( .A(n8975), .B(n1928), .C(tmp_39_i_fu_576_p2[2]), .Y(n1865)
         );
  OAI21X1 U2185 ( .A(n8963), .B(n9893), .C(n6960), .Y(n3984) );
  OAI21X1 U2188 ( .A(n8976), .B(n9892), .C(n7433), .Y(n3985) );
  NAND3X1 U2189 ( .A(ap_CS_fsm[1]), .B(n1928), .C(tmp_39_i_fu_576_p2[4]), .Y(
        n1869) );
  NAND3X1 U2191 ( .A(n1934), .B(n1935), .C(n1936), .Y(n1933) );
  NOR3X1 U2192 ( .A(n8028), .B(n8026), .C(n8027), .Y(n1936) );
  NAND3X1 U2195 ( .A(tmp_39_i_fu_576_p2[4]), .B(tmp_39_i_fu_576_p2[2]), .C(
        n8253), .Y(n1937) );
  NOR3X1 U2197 ( .A(n6940), .B(p_tmp_i_fu_587_p3[1]), .C(p_tmp_i_fu_587_p3[19]), .Y(n1935) );
  NOR3X1 U2199 ( .A(n7086), .B(p_tmp_i_fu_587_p3[16]), .C(
        p_tmp_i_fu_587_p3[15]), .Y(n1934) );
  NAND3X1 U2201 ( .A(n1943), .B(n1944), .C(n1945), .Y(n1932) );
  NOR3X1 U2202 ( .A(n8291), .B(n1947), .C(n8290), .Y(n1945) );
  NAND3X1 U2205 ( .A(n9884), .B(n9883), .C(n8017), .Y(n1946) );
  NOR3X1 U2207 ( .A(n7800), .B(p_tmp_i_fu_587_p3[27]), .C(
        p_tmp_i_fu_587_p3[26]), .Y(n1944) );
  NOR3X1 U2209 ( .A(n7243), .B(p_tmp_i_fu_587_p3[23]), .C(
        p_tmp_i_fu_587_p3[22]), .Y(n1943) );
  OAI21X1 U2212 ( .A(n8980), .B(n8659), .C(n7662), .Y(n3986) );
  OAI21X1 U2215 ( .A(n8979), .B(n9860), .C(n6579), .Y(n3987) );
  OAI21X1 U2218 ( .A(n8978), .B(n9861), .C(n6261), .Y(n3988) );
  OAI21X1 U2221 ( .A(n8979), .B(n9862), .C(n7456), .Y(n3989) );
  OAI21X1 U2224 ( .A(n8977), .B(n9863), .C(n7276), .Y(n3990) );
  OAI21X1 U2227 ( .A(n8980), .B(n9864), .C(n7110), .Y(n3991) );
  OAI21X1 U2230 ( .A(n8979), .B(n9865), .C(n6959), .Y(n3992) );
  OAI21X1 U2233 ( .A(n8978), .B(n9866), .C(n6821), .Y(n3993) );
  OAI21X1 U2236 ( .A(n8978), .B(n9867), .C(n6466), .Y(n3994) );
  OAI21X1 U2239 ( .A(n8977), .B(n9868), .C(n6173), .Y(n3995) );
  OAI21X1 U2242 ( .A(n8978), .B(n9869), .C(n6172), .Y(n3996) );
  OAI21X1 U2245 ( .A(n8978), .B(n9870), .C(n6100), .Y(n3997) );
  OAI21X1 U2248 ( .A(n8978), .B(n9871), .C(n6040), .Y(n3998) );
  OAI21X1 U2251 ( .A(n8978), .B(n9872), .C(n5056), .Y(n3999) );
  OAI21X1 U2254 ( .A(n8978), .B(n9873), .C(n7455), .Y(n4000) );
  OAI21X1 U2257 ( .A(n8978), .B(n9874), .C(n7275), .Y(n4001) );
  OAI21X1 U2260 ( .A(n8978), .B(n9875), .C(n7109), .Y(n4002) );
  OAI21X1 U2263 ( .A(n8978), .B(n9876), .C(n6958), .Y(n4003) );
  OAI21X1 U2266 ( .A(n8977), .B(n9877), .C(n6260), .Y(n4004) );
  OAI21X1 U2269 ( .A(n8980), .B(n9878), .C(n6099), .Y(n4005) );
  OAI21X1 U2272 ( .A(n8978), .B(n9879), .C(n5055), .Y(n4006) );
  OAI21X1 U2275 ( .A(n8979), .B(n9880), .C(n6357), .Y(n4007) );
  OAI21X1 U2278 ( .A(n8978), .B(n9881), .C(n6039), .Y(n4008) );
  OAI21X1 U2281 ( .A(n8978), .B(n9882), .C(n6820), .Y(n4009) );
  OAI21X1 U2284 ( .A(n8980), .B(n9883), .C(n6171), .Y(n4010) );
  OAI21X1 U2287 ( .A(n8977), .B(n9884), .C(n5054), .Y(n4011) );
  OAI21X1 U2290 ( .A(n8978), .B(n9885), .C(n6465), .Y(n4012) );
  OAI21X1 U2293 ( .A(n8964), .B(n9891), .C(n6356), .Y(n4013) );
  OAI21X1 U2296 ( .A(n8975), .B(n9890), .C(n7257), .Y(n4014) );
  OAI21X1 U2299 ( .A(n8963), .B(n9889), .C(n6819), .Y(n4015) );
  OAI21X1 U2302 ( .A(ap_CS_fsm[1]), .B(n9888), .C(n7093), .Y(n4016) );
  OAI21X1 U2305 ( .A(n8963), .B(n9887), .C(n6694), .Y(n4017) );
  OAI21X1 U2308 ( .A(n8975), .B(n9886), .C(n6943), .Y(n4018) );
  OAI21X1 U2311 ( .A(n8975), .B(n9859), .C(n6347), .Y(n4019) );
  OAI21X1 U2313 ( .A(n8976), .B(n9858), .C(n8302), .Y(n4020) );
  OAI21X1 U2315 ( .A(ap_CS_fsm[1]), .B(n9857), .C(n8059), .Y(n4021) );
  OAI21X1 U2317 ( .A(ap_CS_fsm[1]), .B(n9856), .C(n7837), .Y(n4022) );
  OAI21X1 U2319 ( .A(ap_CS_fsm[1]), .B(n9855), .C(n7624), .Y(n4023) );
  OAI21X1 U2321 ( .A(n8975), .B(n9854), .C(n8301), .Y(n4024) );
  OAI21X1 U2324 ( .A(n8976), .B(n9853), .C(n8058), .Y(n4025) );
  OAI21X1 U2327 ( .A(n8976), .B(n9852), .C(n7836), .Y(n4026) );
  OAI21X1 U2329 ( .A(n8976), .B(n9851), .C(n7623), .Y(n4027) );
  OAI21X1 U2331 ( .A(n8975), .B(n9850), .C(n7432), .Y(n4028) );
  OAI21X1 U2334 ( .A(n8975), .B(n9849), .C(n7256), .Y(n4029) );
  OAI21X1 U2337 ( .A(ap_CS_fsm[1]), .B(n9848), .C(n7092), .Y(n4030) );
  OAI21X1 U2339 ( .A(n8976), .B(n9847), .C(n6942), .Y(n4031) );
  OAI21X1 U2341 ( .A(ap_CS_fsm[1]), .B(n9846), .C(n6809), .Y(n4032) );
  OAI21X1 U2344 ( .A(n8975), .B(n9845), .C(n6685), .Y(n4033) );
  OAI21X1 U2346 ( .A(ap_CS_fsm[1]), .B(n9844), .C(n6570), .Y(n4034) );
  OAI21X1 U2348 ( .A(n8976), .B(n9843), .C(n6457), .Y(n4035) );
  OAI21X1 U2351 ( .A(n8976), .B(n9842), .C(n6348), .Y(n4036) );
  OAI21X1 U2354 ( .A(n8975), .B(n9841), .C(n8300), .Y(n4037) );
  OAI21X1 U2356 ( .A(ap_CS_fsm[1]), .B(n9840), .C(n8057), .Y(n4038) );
  OAI21X1 U2358 ( .A(n8976), .B(n9839), .C(n7835), .Y(n4039) );
  OAI21X1 U2360 ( .A(n8976), .B(n9838), .C(n7622), .Y(n4040) );
  OAI21X1 U2362 ( .A(n8976), .B(n9837), .C(n7431), .Y(n4041) );
  OAI21X1 U2365 ( .A(n8976), .B(n9836), .C(n7255), .Y(n4042) );
  OAI21X1 U2368 ( .A(n8976), .B(n9835), .C(n7091), .Y(n4043) );
  OAI21X1 U2370 ( .A(n8976), .B(n9834), .C(n6941), .Y(n4044) );
  OAI21X1 U2372 ( .A(n8976), .B(n9833), .C(n6808), .Y(n4045) );
  OAI21X1 U2374 ( .A(n8976), .B(n9832), .C(n8060), .Y(n4046) );
  OAI21X1 U2378 ( .A(n8976), .B(n9831), .C(n6684), .Y(n4047) );
  OAI21X1 U2380 ( .A(n8976), .B(n9830), .C(n7838), .Y(n4048) );
  OAI21X1 U2381 ( .A(n8976), .B(n9829), .C(n7838), .Y(n4049) );
  OAI21X1 U2385 ( .A(ap_CS_fsm[1]), .B(n9828), .C(n6569), .Y(n4050) );
  OAI21X1 U2386 ( .A(n8976), .B(n9827), .C(n6569), .Y(n4051) );
  OAI21X1 U2389 ( .A(ap_CS_fsm[1]), .B(n9826), .C(n6456), .Y(n4052) );
  OAI21X1 U2392 ( .A(n8975), .B(n9825), .C(n6347), .Y(n4053) );
  NAND3X1 U2396 ( .A(n2030), .B(n2031), .C(n2032), .Y(n2029) );
  NOR3X1 U2397 ( .A(n7615), .B(n7613), .C(n7614), .Y(n2032) );
  NAND3X1 U2404 ( .A(recentdatapoints_len[4]), .B(recentdatapoints_len[2]), 
        .C(n8016), .Y(n2033) );
  NOR3X1 U2406 ( .A(n7090), .B(recentdatapoints_len[1]), .C(
        recentdatapoints_len[19]), .Y(n2031) );
  NOR3X1 U2410 ( .A(n6939), .B(recentdatapoints_len[16]), .C(
        recentdatapoints_len[15]), .Y(n2030) );
  NAND3X1 U2414 ( .A(n2039), .B(n2040), .C(n2041), .Y(n2028) );
  NOR3X1 U2415 ( .A(n7421), .B(n7419), .C(n7420), .Y(n2041) );
  NAND3X1 U2422 ( .A(n9834), .B(n9835), .C(n8015), .Y(n2042) );
  NOR3X1 U2426 ( .A(n6807), .B(recentdatapoints_len[27]), .C(
        recentdatapoints_len[26]), .Y(n2040) );
  NOR3X1 U2430 ( .A(n7245), .B(recentdatapoints_len[23]), .C(
        recentdatapoints_len[22]), .Y(n2039) );
  NAND3X1 U2436 ( .A(\not_tmp_i_i2_reg_1745[0] ), .B(ap_CS_fsm[11]), .C(
        \recentABools_data_q1[0] ), .Y(n2049) );
  NAND3X1 U2501 ( .A(n2053), .B(n2054), .C(n2055), .Y(n2052) );
  NOR3X1 U2502 ( .A(n7818), .B(n7816), .C(n7817), .Y(n2055) );
  NAND3X1 U2509 ( .A(n9912), .B(n9911), .C(n8258), .Y(n2056) );
  NOR3X1 U2513 ( .A(n7418), .B(tmp_38_i_reg_1550[14]), .C(
        tmp_38_i_reg_1550[13]), .Y(n2054) );
  NOR3X1 U2517 ( .A(n7239), .B(tmp_38_i_reg_1550[10]), .C(tmp_38_i_reg_1550[0]), .Y(n2053) );
  NAND3X1 U2521 ( .A(n2062), .B(n2063), .C(n2064), .Y(n2051) );
  NOR3X1 U2522 ( .A(n8031), .B(n8029), .C(n8030), .Y(n2064) );
  NAND3X1 U2529 ( .A(n9926), .B(n9925), .C(n8259), .Y(n2065) );
  NOR3X1 U2533 ( .A(n8285), .B(tmp_38_i_reg_1550[29]), .C(
        tmp_38_i_reg_1550[28]), .Y(n2063) );
  NOR3X1 U2537 ( .A(n7605), .B(tmp_38_i_reg_1550[25]), .C(
        tmp_38_i_reg_1550[24]), .Y(n2062) );
  AOI22X1 U2544 ( .A(data_read_reg_1495[0]), .B(n8969), .C(data[0]), .D(n8963), 
        .Y(n2071) );
  AOI22X1 U2546 ( .A(data_read_reg_1495[1]), .B(n8968), .C(data[1]), .D(n8658), 
        .Y(n2073) );
  AOI22X1 U2548 ( .A(data_read_reg_1495[2]), .B(n8971), .C(data[2]), .D(n8658), 
        .Y(n2074) );
  AOI22X1 U2550 ( .A(data_read_reg_1495[3]), .B(n8969), .C(data[3]), .D(n8967), 
        .Y(n2075) );
  AOI22X1 U2552 ( .A(data_read_reg_1495[4]), .B(n8968), .C(data[4]), .D(n8658), 
        .Y(n2076) );
  AOI22X1 U2554 ( .A(data_read_reg_1495[5]), .B(n8971), .C(data[5]), .D(n8658), 
        .Y(n2077) );
  AOI22X1 U2556 ( .A(data_read_reg_1495[6]), .B(n8970), .C(data[6]), .D(n8658), 
        .Y(n2078) );
  AOI22X1 U2558 ( .A(data_read_reg_1495[7]), .B(n8968), .C(data[7]), .D(n8658), 
        .Y(n2079) );
  AOI22X1 U2560 ( .A(data_read_reg_1495[8]), .B(n8968), .C(data[8]), .D(n8658), 
        .Y(n2080) );
  AOI22X1 U2562 ( .A(data_read_reg_1495[9]), .B(n8968), .C(data[9]), .D(n8658), 
        .Y(n2081) );
  AOI22X1 U2564 ( .A(data_read_reg_1495[10]), .B(n8968), .C(data[10]), .D(
        n8967), .Y(n2082) );
  AOI22X1 U2566 ( .A(data_read_reg_1495[11]), .B(n8968), .C(data[11]), .D(
        n8658), .Y(n2083) );
  AOI22X1 U2568 ( .A(data_read_reg_1495[12]), .B(n8968), .C(data[12]), .D(
        n8967), .Y(n2084) );
  AOI22X1 U2570 ( .A(data_read_reg_1495[13]), .B(n8968), .C(data[13]), .D(
        n8658), .Y(n2085) );
  AOI22X1 U2572 ( .A(data_read_reg_1495[14]), .B(n8968), .C(data[14]), .D(
        n8967), .Y(n2086) );
  AOI22X1 U2574 ( .A(data_read_reg_1495[15]), .B(n8968), .C(data[15]), .D(
        n8658), .Y(n2087) );
  AOI22X1 U2576 ( .A(vthresh[0]), .B(n8940), .C(v_thresh[0]), .D(n8956), .Y(
        n2088) );
  AOI22X1 U2578 ( .A(vthresh[1]), .B(n8940), .C(v_thresh[1]), .D(n8956), .Y(
        n2091) );
  AOI22X1 U2580 ( .A(vthresh[2]), .B(n8945), .C(v_thresh[2]), .D(n8960), .Y(
        n2092) );
  AOI22X1 U2582 ( .A(vthresh[3]), .B(n8945), .C(v_thresh[3]), .D(n8960), .Y(
        n2093) );
  AOI22X1 U2584 ( .A(vthresh[4]), .B(n8945), .C(v_thresh[4]), .D(n8960), .Y(
        n2094) );
  AOI22X1 U2586 ( .A(vthresh[5]), .B(n8944), .C(v_thresh[5]), .D(n8960), .Y(
        n2095) );
  AOI22X1 U2588 ( .A(vthresh[6]), .B(n8944), .C(v_thresh[6]), .D(n8960), .Y(
        n2096) );
  AOI22X1 U2590 ( .A(vthresh[7]), .B(n8944), .C(v_thresh[7]), .D(n8960), .Y(
        n2097) );
  AOI22X1 U2592 ( .A(vthresh[8]), .B(n8944), .C(v_thresh[8]), .D(n8960), .Y(
        n2098) );
  AOI22X1 U2594 ( .A(vthresh[9]), .B(n8944), .C(v_thresh[9]), .D(n8960), .Y(
        n2099) );
  AOI22X1 U2596 ( .A(vthresh[10]), .B(n8944), .C(v_thresh[10]), .D(n8960), .Y(
        n2100) );
  AOI22X1 U2598 ( .A(vthresh[11]), .B(n8944), .C(v_thresh[11]), .D(n8960), .Y(
        n2101) );
  AOI22X1 U2600 ( .A(vthresh[12]), .B(n8944), .C(v_thresh[12]), .D(n8960), .Y(
        n2102) );
  AOI22X1 U2602 ( .A(vthresh[13]), .B(n8944), .C(v_thresh[13]), .D(n8959), .Y(
        n2103) );
  AOI22X1 U2604 ( .A(vthresh[14]), .B(n8944), .C(v_thresh[14]), .D(n8959), .Y(
        n2104) );
  AOI22X1 U2606 ( .A(vthresh[15]), .B(n8944), .C(v_thresh[15]), .D(n8959), .Y(
        n2105) );
  AOI22X1 U2608 ( .A(vthresh[16]), .B(n8942), .C(v_thresh[16]), .D(n8959), .Y(
        n2106) );
  AOI22X1 U2610 ( .A(vthresh[17]), .B(n8943), .C(v_thresh[17]), .D(n8959), .Y(
        n2107) );
  AOI22X1 U2612 ( .A(vthresh[18]), .B(n8944), .C(v_thresh[18]), .D(n8959), .Y(
        n2108) );
  AOI22X1 U2614 ( .A(vthresh[19]), .B(n8944), .C(v_thresh[19]), .D(n8959), .Y(
        n2109) );
  AOI22X1 U2616 ( .A(vthresh[20]), .B(n8943), .C(v_thresh[20]), .D(n8959), .Y(
        n2110) );
  AOI22X1 U2618 ( .A(vthresh[21]), .B(n8943), .C(v_thresh[21]), .D(n8959), .Y(
        n2111) );
  AOI22X1 U2620 ( .A(vthresh[22]), .B(n8943), .C(v_thresh[22]), .D(n8959), .Y(
        n2112) );
  AOI22X1 U2622 ( .A(vthresh[23]), .B(n8943), .C(v_thresh[23]), .D(n8959), .Y(
        n2113) );
  AOI22X1 U2624 ( .A(vthresh[24]), .B(n8943), .C(v_thresh[24]), .D(n8958), .Y(
        n2114) );
  AOI22X1 U2626 ( .A(vthresh[25]), .B(n8943), .C(v_thresh[25]), .D(n8958), .Y(
        n2115) );
  AOI22X1 U2628 ( .A(vthresh[26]), .B(n8943), .C(v_thresh[26]), .D(n8958), .Y(
        n2116) );
  AOI22X1 U2630 ( .A(vthresh[27]), .B(n8943), .C(v_thresh[27]), .D(n8958), .Y(
        n2117) );
  AOI22X1 U2632 ( .A(vthresh[28]), .B(n8943), .C(v_thresh[28]), .D(n8958), .Y(
        n2118) );
  AOI22X1 U2634 ( .A(vthresh[29]), .B(n8943), .C(v_thresh[29]), .D(n8958), .Y(
        n2119) );
  AOI22X1 U2636 ( .A(vthresh[30]), .B(n8943), .C(v_thresh[30]), .D(n8958), .Y(
        n2120) );
  AOI22X1 U2638 ( .A(vthresh[31]), .B(n8943), .C(v_thresh[31]), .D(n8958), .Y(
        n2121) );
  AOI22X1 U2640 ( .A(athresh[0]), .B(n8941), .C(a_thresh[0]), .D(n8958), .Y(
        n2122) );
  AOI22X1 U2642 ( .A(athresh[1]), .B(n8942), .C(a_thresh[1]), .D(n8958), .Y(
        n2123) );
  AOI22X1 U2644 ( .A(athresh[2]), .B(n8942), .C(a_thresh[2]), .D(n8958), .Y(
        n2124) );
  AOI22X1 U2646 ( .A(athresh[3]), .B(n8942), .C(a_thresh[3]), .D(n8957), .Y(
        n2125) );
  AOI22X1 U2648 ( .A(athresh[4]), .B(n8942), .C(a_thresh[4]), .D(n8957), .Y(
        n2126) );
  AOI22X1 U2650 ( .A(athresh[5]), .B(n8942), .C(a_thresh[5]), .D(n8957), .Y(
        n2127) );
  AOI22X1 U2652 ( .A(athresh[6]), .B(n8942), .C(a_thresh[6]), .D(n8957), .Y(
        n2128) );
  AOI22X1 U2654 ( .A(athresh[7]), .B(n8942), .C(a_thresh[7]), .D(n8957), .Y(
        n2129) );
  AOI22X1 U2656 ( .A(athresh[8]), .B(n8942), .C(a_thresh[8]), .D(n8957), .Y(
        n2130) );
  AOI22X1 U2658 ( .A(athresh[9]), .B(n8942), .C(a_thresh[9]), .D(n8957), .Y(
        n2131) );
  AOI22X1 U2660 ( .A(athresh[10]), .B(n8942), .C(a_thresh[10]), .D(n8957), .Y(
        n2132) );
  AOI22X1 U2662 ( .A(athresh[11]), .B(n8942), .C(a_thresh[11]), .D(n8957), .Y(
        n2133) );
  AOI22X1 U2664 ( .A(athresh[12]), .B(n8941), .C(a_thresh[12]), .D(n8957), .Y(
        n2134) );
  AOI22X1 U2666 ( .A(athresh[13]), .B(n8942), .C(a_thresh[13]), .D(n8957), .Y(
        n2135) );
  AOI22X1 U2668 ( .A(athresh[14]), .B(n8941), .C(a_thresh[14]), .D(n8956), .Y(
        n2136) );
  AOI22X1 U2670 ( .A(athresh[15]), .B(n8941), .C(a_thresh[15]), .D(n8956), .Y(
        n2137) );
  AOI22X1 U2672 ( .A(athresh[16]), .B(n8940), .C(a_thresh[16]), .D(n8956), .Y(
        n2138) );
  AOI22X1 U2674 ( .A(athresh[17]), .B(n8941), .C(a_thresh[17]), .D(n8956), .Y(
        n2139) );
  AOI22X1 U2676 ( .A(athresh[18]), .B(n8941), .C(a_thresh[18]), .D(n8956), .Y(
        n2140) );
  AOI22X1 U2678 ( .A(athresh[19]), .B(n8941), .C(a_thresh[19]), .D(n8956), .Y(
        n2141) );
  AOI22X1 U2680 ( .A(athresh[20]), .B(n8941), .C(a_thresh[20]), .D(n8956), .Y(
        n2142) );
  AOI22X1 U2682 ( .A(athresh[21]), .B(n8941), .C(a_thresh[21]), .D(n8956), .Y(
        n2143) );
  AOI22X1 U2684 ( .A(athresh[22]), .B(n8941), .C(a_thresh[22]), .D(n8956), .Y(
        n2144) );
  AOI22X1 U2686 ( .A(athresh[23]), .B(n8941), .C(a_thresh[23]), .D(n8956), .Y(
        n2145) );
  AOI22X1 U2688 ( .A(athresh[24]), .B(n8940), .C(a_thresh[24]), .D(n8956), .Y(
        n2146) );
  AOI22X1 U2690 ( .A(athresh[25]), .B(n8941), .C(a_thresh[25]), .D(n8958), .Y(
        n2147) );
  AOI22X1 U2692 ( .A(athresh[26]), .B(n8941), .C(a_thresh[26]), .D(n8960), .Y(
        n2148) );
  AOI22X1 U2694 ( .A(athresh[27]), .B(n8940), .C(a_thresh[27]), .D(n8958), .Y(
        n2149) );
  AOI22X1 U2696 ( .A(athresh[28]), .B(n8940), .C(a_thresh[28]), .D(n8959), .Y(
        n2150) );
  AOI22X1 U2698 ( .A(athresh[29]), .B(n8940), .C(a_thresh[29]), .D(n8957), .Y(
        n2151) );
  AOI22X1 U2700 ( .A(athresh[30]), .B(n8940), .C(a_thresh[30]), .D(n8957), .Y(
        n2152) );
  AOI22X1 U2702 ( .A(athresh[31]), .B(n8940), .C(a_thresh[31]), .D(n8957), .Y(
        n2153) );
  OAI21X1 U2704 ( .A(ap_CS_fsm[12]), .B(n9385), .C(n8303), .Y(n4168) );
  OAI21X1 U2706 ( .A(n10366), .B(n2156), .C(n6055), .Y(n4169) );
  OAI21X1 U2709 ( .A(n10369), .B(n2156), .C(n6194), .Y(n4170) );
  OAI21X1 U2712 ( .A(n10371), .B(n2156), .C(n6284), .Y(n4171) );
  OAI21X1 U2715 ( .A(n10374), .B(n2156), .C(n6385), .Y(n4172) );
  OAI21X1 U2718 ( .A(n10376), .B(n2156), .C(n6490), .Y(n4173) );
  OAI21X1 U2721 ( .A(n10378), .B(n2156), .C(n6602), .Y(n4174) );
  OAI21X1 U2724 ( .A(n10380), .B(n2156), .C(n6719), .Y(n4175) );
  OAI21X1 U2727 ( .A(n10383), .B(n2156), .C(n6846), .Y(n4176) );
  OAI21X1 U2730 ( .A(n10385), .B(n2156), .C(n6120), .Y(n4177) );
  OAI21X1 U2733 ( .A(n10389), .B(n2156), .C(n6987), .Y(n4178) );
  OAI21X1 U2736 ( .A(n10391), .B(n2156), .C(n7479), .Y(n4179) );
  OAI21X1 U2739 ( .A(n10395), .B(n2156), .C(n7683), .Y(n4180) );
  OAI21X1 U2742 ( .A(n10397), .B(n2156), .C(n7136), .Y(n4181) );
  OAI21X1 U2745 ( .A(n10400), .B(n2156), .C(n7300), .Y(n4182) );
  OAI21X1 U2748 ( .A(n10402), .B(n2156), .C(n8150), .Y(n4183) );
  OAI21X1 U2751 ( .A(n10406), .B(n2156), .C(n6195), .Y(n4184) );
  OAI21X1 U2754 ( .A(n10408), .B(n2156), .C(n6286), .Y(n4185) );
  OAI21X1 U2757 ( .A(n10410), .B(n2156), .C(n6387), .Y(n4186) );
  OAI21X1 U2760 ( .A(n10412), .B(n2156), .C(n6494), .Y(n4187) );
  OAI21X1 U2763 ( .A(n10416), .B(n2156), .C(n6606), .Y(n4188) );
  OAI21X1 U2766 ( .A(n10418), .B(n2156), .C(n6723), .Y(n4189) );
  OAI21X1 U2769 ( .A(n10421), .B(n2156), .C(n7482), .Y(n4190) );
  OAI21X1 U2772 ( .A(n10423), .B(n2156), .C(n7686), .Y(n4191) );
  OAI21X1 U2775 ( .A(n10427), .B(n2156), .C(n7901), .Y(n4192) );
  OAI21X1 U2778 ( .A(n10429), .B(n2156), .C(n6850), .Y(n4193) );
  OAI21X1 U2781 ( .A(n10432), .B(n2156), .C(n6990), .Y(n4194) );
  OAI21X1 U2784 ( .A(n10434), .B(n2156), .C(n7139), .Y(n4195) );
  OAI21X1 U2787 ( .A(n10438), .B(n2156), .C(n7303), .Y(n4196) );
  OAI21X1 U2790 ( .A(n10440), .B(n2156), .C(n8152), .Y(n4197) );
  OAI21X1 U2793 ( .A(n10442), .B(n2156), .C(n7484), .Y(n4198) );
  OAI21X1 U2796 ( .A(n10444), .B(n2156), .C(n7687), .Y(n4199) );
  OAI21X1 U2799 ( .A(n10448), .B(n2156), .C(n7903), .Y(n4200) );
  OAI21X1 U2801 ( .A(N495), .B(n10240), .C(ap_CS_fsm[7]), .Y(n2156) );
  NAND3X1 U2804 ( .A(n10674), .B(N503), .C(\tmp_25_reg_1777[0] ), .Y(n585) );
  AOI22X1 U2808 ( .A(i_11_fu_1179_p2[4]), .B(n10279), .C(i_12_fu_1191_p2[4]), 
        .D(i_11_fu_1179_p2[31]), .Y(n2190) );
  AOI22X1 U2810 ( .A(i_11_fu_1179_p2[3]), .B(n10279), .C(i_12_fu_1191_p2[3]), 
        .D(i_11_fu_1179_p2[31]), .Y(n2192) );
  AOI22X1 U2812 ( .A(i_11_fu_1179_p2[2]), .B(n10279), .C(i_12_fu_1191_p2[2]), 
        .D(i_11_fu_1179_p2[31]), .Y(n2193) );
  AOI22X1 U2814 ( .A(i_11_fu_1179_p2[1]), .B(n10279), .C(n10305), .D(
        i_11_fu_1179_p2[31]), .Y(n2194) );
  AOI22X1 U2816 ( .A(i_12_fu_1191_p2[0]), .B(n10279), .C(i_12_fu_1191_p2[0]), 
        .D(i_11_fu_1179_p2[31]), .Y(n2195) );
  AOI22X1 U2819 ( .A(i_5_fu_854_p2[4]), .B(n9997), .C(i_6_fu_866_p2[4]), .D(
        i_5_fu_854_p2[31]), .Y(n2196) );
  AOI22X1 U2821 ( .A(i_5_fu_854_p2[3]), .B(n9997), .C(i_6_fu_866_p2[3]), .D(
        i_5_fu_854_p2[31]), .Y(n2198) );
  AOI22X1 U2823 ( .A(i_5_fu_854_p2[2]), .B(n9997), .C(i_6_fu_866_p2[2]), .D(
        i_5_fu_854_p2[31]), .Y(n2199) );
  AOI22X1 U2825 ( .A(i_5_fu_854_p2[1]), .B(n9997), .C(n10023), .D(
        i_5_fu_854_p2[31]), .Y(n2200) );
  AOI22X1 U2827 ( .A(i_6_fu_866_p2[0]), .B(n9997), .C(i_6_fu_866_p2[0]), .D(
        i_5_fu_854_p2[31]), .Y(n2201) );
  OAI21X1 U2829 ( .A(n10738), .B(n2202), .C(n8172), .Y(n4214) );
  OAI21X1 U2832 ( .A(n10736), .B(n2202), .C(n7926), .Y(n4215) );
  OAI21X1 U2835 ( .A(n10734), .B(n2202), .C(n7710), .Y(n4216) );
  OAI21X1 U2838 ( .A(n10732), .B(n2202), .C(n7510), .Y(n4217) );
  OAI21X1 U2841 ( .A(n10730), .B(n2202), .C(n7330), .Y(n4218) );
  OAI21X1 U2844 ( .A(n10728), .B(n2202), .C(n7166), .Y(n4219) );
  OAI21X1 U2847 ( .A(n10726), .B(n2202), .C(n7015), .Y(n4220) );
  OAI21X1 U2850 ( .A(n10724), .B(n2202), .C(n6875), .Y(n4221) );
  OAI21X1 U2853 ( .A(n10722), .B(n2202), .C(n6748), .Y(n4222) );
  OAI21X1 U2856 ( .A(n10720), .B(n2202), .C(n6628), .Y(n4223) );
  OAI21X1 U2859 ( .A(n10718), .B(n2202), .C(n6516), .Y(n4224) );
  OAI21X1 U2862 ( .A(n10716), .B(n2202), .C(n6407), .Y(n4225) );
  OAI21X1 U2865 ( .A(n10714), .B(n2202), .C(n7924), .Y(n4226) );
  OAI21X1 U2868 ( .A(n10712), .B(n2202), .C(n7707), .Y(n4227) );
  OAI21X1 U2871 ( .A(n10710), .B(n2202), .C(n7507), .Y(n4228) );
  OAI21X1 U2874 ( .A(n10708), .B(n2202), .C(n7328), .Y(n4229) );
  OAI21X1 U2877 ( .A(n10706), .B(n2202), .C(n7163), .Y(n4230) );
  OAI21X1 U2880 ( .A(n10704), .B(n2202), .C(n6298), .Y(n4231) );
  OAI21X1 U2883 ( .A(n10702), .B(n2202), .C(n6206), .Y(n4232) );
  OAI21X1 U2886 ( .A(n10700), .B(n2202), .C(n6126), .Y(n4233) );
  OAI21X1 U2889 ( .A(n10698), .B(n2202), .C(n7013), .Y(n4234) );
  OAI21X1 U2892 ( .A(n10696), .B(n2202), .C(n8169), .Y(n4235) );
  OAI21X1 U2895 ( .A(n10694), .B(n2202), .C(n6872), .Y(n4236) );
  OAI21X1 U2898 ( .A(n10692), .B(n2202), .C(n6745), .Y(n4237) );
  OAI21X1 U2901 ( .A(n10690), .B(n2202), .C(n7923), .Y(n4238) );
  OAI21X1 U2904 ( .A(n10687), .B(n2202), .C(n7505), .Y(n4239) );
  OAI21X1 U2907 ( .A(n10684), .B(n2202), .C(n7705), .Y(n4240) );
  OAI21X1 U2910 ( .A(n10682), .B(n2202), .C(n7326), .Y(n4241) );
  OAI21X1 U2913 ( .A(n10680), .B(n2202), .C(n7160), .Y(n4242) );
  OAI21X1 U2916 ( .A(n10678), .B(n2202), .C(n6625), .Y(n4243) );
  OAI21X1 U2919 ( .A(n10672), .B(n2202), .C(n6512), .Y(n4244) );
  OAI21X1 U2922 ( .A(ap_CS_fsm[12]), .B(n10810), .C(n8303), .Y(n4245) );
  OAI21X1 U2926 ( .A(n7260), .B(n8934), .C(n4819), .Y(n4246) );
  AOI22X1 U2927 ( .A(recentABools_len_new_reg_385[30]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[30]), .D(n2403), .Y(n2240)
         );
  OAI21X1 U2928 ( .A(n6166), .B(n8934), .C(n4818), .Y(n4247) );
  AOI22X1 U2929 ( .A(recentABools_len_new_reg_385[29]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[29]), .D(n2403), .Y(n2244)
         );
  OAI21X1 U2930 ( .A(n6688), .B(n8934), .C(n4817), .Y(n4248) );
  AOI22X1 U2931 ( .A(recentABools_len_new_reg_385[28]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[28]), .D(n2403), .Y(n2246)
         );
  OAI21X1 U2932 ( .A(n7646), .B(n8934), .C(n7323), .Y(n4249) );
  AOI22X1 U2933 ( .A(recentABools_len_new_reg_385[27]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[27]), .D(n2403), .Y(n2248)
         );
  OAI21X1 U2934 ( .A(n6813), .B(n8934), .C(n4816), .Y(n4250) );
  AOI22X1 U2935 ( .A(recentABools_len_new_reg_385[26]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[26]), .D(n2403), .Y(n2250)
         );
  OAI21X1 U2936 ( .A(n6948), .B(n8934), .C(n4815), .Y(n4251) );
  AOI22X1 U2937 ( .A(recentABools_len_new_reg_385[25]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[25]), .D(n2403), .Y(n2252)
         );
  OAI21X1 U2938 ( .A(n6573), .B(n2239), .C(n4814), .Y(n4252) );
  AOI22X1 U2939 ( .A(recentABools_len_new_reg_385[24]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[24]), .D(n2403), .Y(n2254)
         );
  OAI21X1 U2940 ( .A(n8401), .B(n8934), .C(n7159), .Y(n4253) );
  AOI22X1 U2941 ( .A(recentABools_len_new_reg_385[23]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[23]), .D(n2403), .Y(n2256)
         );
  OAI21X1 U2942 ( .A(n7100), .B(n2239), .C(n4813), .Y(n4254) );
  AOI22X1 U2943 ( .A(recentABools_len_new_reg_385[22]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[22]), .D(n2403), .Y(n2258)
         );
  OAI21X1 U2944 ( .A(n7265), .B(n8934), .C(n4812), .Y(n4255) );
  AOI22X1 U2945 ( .A(recentABools_len_new_reg_385[21]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[21]), .D(n2403), .Y(n2260)
         );
  OAI21X1 U2946 ( .A(n6460), .B(n2239), .C(n4811), .Y(n4256) );
  AOI22X1 U2947 ( .A(recentABools_len_new_reg_385[20]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[20]), .D(n2403), .Y(n2262)
         );
  OAI21X1 U2948 ( .A(n7864), .B(n8934), .C(n7500), .Y(n4257) );
  AOI22X1 U2949 ( .A(recentABools_len_new_reg_385[19]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[19]), .D(n2403), .Y(n2264)
         );
  OAI21X1 U2950 ( .A(n7443), .B(n8934), .C(n4810), .Y(n4258) );
  AOI22X1 U2951 ( .A(recentABools_len_new_reg_385[18]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[18]), .D(n2403), .Y(n2266)
         );
  OAI21X1 U2952 ( .A(n6351), .B(n2239), .C(n4809), .Y(n4259) );
  AOI22X1 U2953 ( .A(recentABools_len_new_reg_385[17]), .B(n8932), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[17]), .D(n8890), .Y(n2268)
         );
  OAI21X1 U2954 ( .A(n6254), .B(n2239), .C(n4808), .Y(n4260) );
  AOI22X1 U2955 ( .A(recentABools_len_new_reg_385[16]), .B(n8932), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[16]), .D(n2403), .Y(n2270)
         );
  OAI21X1 U2956 ( .A(n8114), .B(n8934), .C(n7321), .Y(n4261) );
  AOI22X1 U2957 ( .A(recentABools_len_new_reg_385[15]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[15]), .D(n8890), .Y(n2272)
         );
  OAI21X1 U2958 ( .A(n8103), .B(n8934), .C(n7008), .Y(n4262) );
  AOI22X1 U2959 ( .A(recentABools_len_new_reg_385[14]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[14]), .D(n2403), .Y(n2274)
         );
  OAI21X1 U2960 ( .A(n7642), .B(n2239), .C(n4807), .Y(n4263) );
  AOI22X1 U2961 ( .A(recentABools_len_new_reg_385[13]), .B(n8932), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[13]), .D(n8890), .Y(n2276)
         );
  OAI21X1 U2962 ( .A(n7439), .B(n8934), .C(n4806), .Y(n4264) );
  AOI22X1 U2963 ( .A(recentABools_len_new_reg_385[12]), .B(n8932), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[12]), .D(n2403), .Y(n2278)
         );
  OAI21X1 U2964 ( .A(n8399), .B(n8934), .C(n7157), .Y(n4265) );
  AOI22X1 U2965 ( .A(recentABools_len_new_reg_385[11]), .B(n8932), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[11]), .D(n8890), .Y(n2280)
         );
  OAI21X1 U2966 ( .A(n7860), .B(n8934), .C(n7498), .Y(n4266) );
  AOI22X1 U2967 ( .A(recentABools_len_new_reg_385[10]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[10]), .D(n2403), .Y(n2282)
         );
  OAI21X1 U2968 ( .A(n7862), .B(n2239), .C(n6867), .Y(n4267) );
  AOI22X1 U2969 ( .A(recentABools_len_new_reg_385[9]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[9]), .D(n8890), .Y(n2284)
         );
  OAI21X1 U2970 ( .A(n8407), .B(n8934), .C(n6739), .Y(n4268) );
  AOI22X1 U2971 ( .A(recentABools_len_new_reg_385[8]), .B(n8932), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[8]), .D(n2403), .Y(n2286)
         );
  OAI21X1 U2972 ( .A(n8112), .B(n8934), .C(n6621), .Y(n4269) );
  AOI22X1 U2973 ( .A(recentABools_len_new_reg_385[7]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[7]), .D(n8890), .Y(n2288)
         );
  OAI21X1 U2974 ( .A(n7644), .B(n2239), .C(n6509), .Y(n4270) );
  AOI22X1 U2975 ( .A(recentABools_len_new_reg_385[6]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[6]), .D(n8890), .Y(n2290)
         );
  OAI21X1 U2976 ( .A(n7441), .B(n2239), .C(n6402), .Y(n4271) );
  AOI22X1 U2977 ( .A(recentABools_len_new_reg_385[5]), .B(n8932), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[5]), .D(n8890), .Y(n2292)
         );
  OAI21X1 U2978 ( .A(n10536), .B(n8934), .C(n7319), .Y(n4272) );
  AOI22X1 U2979 ( .A(recentABools_len_new_reg_385[4]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[4]), .D(n8890), .Y(n2294)
         );
  OAI21X1 U2981 ( .A(n10537), .B(n8934), .C(n7006), .Y(n4273) );
  AOI22X1 U2982 ( .A(recentABools_len_new_reg_385[3]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[3]), .D(n8890), .Y(n2296)
         );
  OAI21X1 U2984 ( .A(n10538), .B(n2239), .C(n6296), .Y(n4274) );
  AOI22X1 U2985 ( .A(recentABools_len_new_reg_385[2]), .B(n8932), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[2]), .D(n8890), .Y(n2298)
         );
  OAI21X1 U2987 ( .A(n10539), .B(n8934), .C(n7497), .Y(n4275) );
  AOI22X1 U2988 ( .A(recentABools_len_new_reg_385[1]), .B(n8932), .C(n10574), 
        .D(n8890), .Y(n2300) );
  OAI21X1 U2990 ( .A(n8392), .B(n2239), .C(n7704), .Y(n4276) );
  AOI22X1 U2991 ( .A(recentABools_len_new_reg_385[0]), .B(n2241), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[0]), .D(n8890), .Y(n2302)
         );
  OAI21X1 U2992 ( .A(n4689), .B(n8934), .C(n7937), .Y(n4277) );
  AOI22X1 U2993 ( .A(n8932), .B(sum_1_reg_376[31]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[31]), .Y(n2303) );
  OAI21X1 U2995 ( .A(n8489), .B(n2239), .C(n6094), .Y(n4278) );
  AOI22X1 U2996 ( .A(n2241), .B(sum_1_reg_376[30]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[30]), .Y(n2304) );
  OAI21X1 U2998 ( .A(n8458), .B(n8934), .C(n7152), .Y(n4279) );
  AOI22X1 U2999 ( .A(n2241), .B(sum_1_reg_376[29]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[29]), .Y(n2305) );
  OAI21X1 U3001 ( .A(n8457), .B(n8934), .C(n6864), .Y(n4280) );
  AOI22X1 U3002 ( .A(n8932), .B(sum_1_reg_376[28]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[28]), .Y(n2306) );
  OAI21X1 U3004 ( .A(n8456), .B(n2239), .C(n6619), .Y(n4281) );
  AOI22X1 U3005 ( .A(n8932), .B(sum_1_reg_376[27]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[27]), .Y(n2307) );
  OAI21X1 U3007 ( .A(n8455), .B(n8934), .C(n6736), .Y(n4282) );
  AOI22X1 U3008 ( .A(n2241), .B(sum_1_reg_376[26]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[26]), .Y(n2308) );
  OAI21X1 U3010 ( .A(n8454), .B(n8934), .C(n7002), .Y(n4283) );
  AOI22X1 U3011 ( .A(n8932), .B(sum_1_reg_376[25]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[25]), .Y(n2309) );
  OAI21X1 U3013 ( .A(n8453), .B(n2239), .C(n7315), .Y(n4284) );
  AOI22X1 U3014 ( .A(n8932), .B(sum_1_reg_376[24]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[24]), .Y(n2310) );
  OAI21X1 U3016 ( .A(n8452), .B(n8934), .C(n6505), .Y(n4285) );
  AOI22X1 U3017 ( .A(n8932), .B(sum_1_reg_376[23]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[23]), .Y(n2311) );
  OAI21X1 U3019 ( .A(n8451), .B(n8934), .C(n7698), .Y(n4286) );
  AOI22X1 U3020 ( .A(n8932), .B(sum_1_reg_376[22]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[22]), .Y(n2312) );
  OAI21X1 U3022 ( .A(n8450), .B(n8934), .C(n7914), .Y(n4287) );
  AOI22X1 U3023 ( .A(n8932), .B(sum_1_reg_376[21]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[21]), .Y(n2313) );
  OAI21X1 U3025 ( .A(n8449), .B(n8934), .C(n7495), .Y(n4288) );
  AOI22X1 U3026 ( .A(n8932), .B(sum_1_reg_376[20]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[20]), .Y(n2314) );
  OAI21X1 U3028 ( .A(n8448), .B(n8934), .C(n6398), .Y(n4289) );
  AOI22X1 U3029 ( .A(n8932), .B(sum_1_reg_376[19]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[19]), .Y(n2315) );
  OAI21X1 U3031 ( .A(n8447), .B(n8934), .C(n6294), .Y(n4290) );
  AOI22X1 U3032 ( .A(n8932), .B(sum_1_reg_376[18]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[18]), .Y(n2316) );
  OAI21X1 U3034 ( .A(n8446), .B(n8934), .C(n6203), .Y(n4291) );
  AOI22X1 U3035 ( .A(n8932), .B(sum_1_reg_376[17]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[17]), .Y(n2317) );
  OAI21X1 U3037 ( .A(n8445), .B(n8934), .C(n6862), .Y(n4292) );
  AOI22X1 U3038 ( .A(n8932), .B(sum_1_reg_376[16]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[16]), .Y(n2318) );
  OAI21X1 U3040 ( .A(n8444), .B(n8934), .C(n7149), .Y(n4293) );
  AOI22X1 U3041 ( .A(n8932), .B(sum_1_reg_376[15]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[15]), .Y(n2319) );
  OAI21X1 U3043 ( .A(n8443), .B(n8934), .C(n6734), .Y(n4294) );
  AOI22X1 U3044 ( .A(n8932), .B(sum_1_reg_376[14]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[14]), .Y(n2320) );
  OAI21X1 U3046 ( .A(n8442), .B(n8934), .C(n6617), .Y(n4295) );
  AOI22X1 U3047 ( .A(n8932), .B(sum_1_reg_376[13]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[13]), .Y(n2321) );
  OAI21X1 U3049 ( .A(n8441), .B(n2239), .C(n6293), .Y(n4296) );
  AOI22X1 U3050 ( .A(n2241), .B(sum_1_reg_376[12]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[12]), .Y(n2322) );
  OAI21X1 U3052 ( .A(n8440), .B(n8934), .C(n7313), .Y(n4297) );
  AOI22X1 U3053 ( .A(n8932), .B(sum_1_reg_376[11]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[11]), .Y(n2323) );
  OAI21X1 U3055 ( .A(n8439), .B(n8934), .C(n7000), .Y(n4298) );
  AOI22X1 U3056 ( .A(n2241), .B(sum_1_reg_376[10]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[10]), .Y(n2324) );
  OAI21X1 U3058 ( .A(n8438), .B(n2239), .C(n7912), .Y(n4299) );
  AOI22X1 U3059 ( .A(n8932), .B(sum_1_reg_376[9]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[9]), .Y(n2325) );
  OAI21X1 U3061 ( .A(n8437), .B(n2239), .C(n7696), .Y(n4300) );
  AOI22X1 U3062 ( .A(n2241), .B(sum_1_reg_376[8]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[8]), .Y(n2326) );
  OAI21X1 U3064 ( .A(n8436), .B(n2239), .C(n7493), .Y(n4301) );
  AOI22X1 U3065 ( .A(n8932), .B(sum_1_reg_376[7]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[7]), .Y(n2327) );
  OAI21X1 U3067 ( .A(n8435), .B(n2239), .C(n6503), .Y(n4302) );
  AOI22X1 U3068 ( .A(n2241), .B(sum_1_reg_376[6]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[6]), .Y(n2328) );
  OAI21X1 U3070 ( .A(n8434), .B(n2239), .C(n6396), .Y(n4303) );
  AOI22X1 U3071 ( .A(n8932), .B(sum_1_reg_376[5]), .C(n2403), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[5]), .Y(n2329) );
  OAI21X1 U3073 ( .A(n8433), .B(n2239), .C(n6201), .Y(n4304) );
  AOI22X1 U3074 ( .A(n2241), .B(sum_1_reg_376[4]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[4]), .Y(n2330) );
  OAI21X1 U3076 ( .A(n8432), .B(n2239), .C(n7148), .Y(n4305) );
  AOI22X1 U3077 ( .A(n8932), .B(sum_1_reg_376[3]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[3]), .Y(n2331) );
  OAI21X1 U3079 ( .A(n8431), .B(n8934), .C(n6859), .Y(n4306) );
  AOI22X1 U3080 ( .A(n2241), .B(sum_1_reg_376[2]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[2]), .Y(n2332) );
  OAI21X1 U3082 ( .A(n8430), .B(n2239), .C(n6731), .Y(n4307) );
  AOI22X1 U3083 ( .A(n8932), .B(sum_1_reg_376[1]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[1]), .Y(n2333) );
  OAI21X1 U3085 ( .A(n8662), .B(n8934), .C(n6614), .Y(n4308) );
  AOI22X1 U3086 ( .A(n2241), .B(sum_1_reg_376[0]), .C(n8890), .D(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[0]), .Y(n2334) );
  OAI21X1 U3088 ( .A(ap_CS_fsm[12]), .B(n10669), .C(n8166), .Y(n4309) );
  AOI22X1 U3089 ( .A(recentABools_len_new_reg_385[31]), .B(n8931), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[31]), .D(n8657), .Y(n2336)
         );
  OAI21X1 U3090 ( .A(ap_CS_fsm[12]), .B(n10573), .C(n7153), .Y(n4310) );
  AOI22X1 U3091 ( .A(n8931), .B(recentABools_len_new_reg_385[30]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[30]), .D(n8657), .Y(n2340)
         );
  OAI21X1 U3092 ( .A(ap_CS_fsm[12]), .B(n10633), .C(n7502), .Y(n4311) );
  AOI22X1 U3093 ( .A(n8931), .B(recentABools_len_new_reg_385[29]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[29]), .D(n8657), .Y(n2342)
         );
  OAI21X1 U3094 ( .A(ap_CS_fsm[12]), .B(n10632), .C(n7324), .Y(n4312) );
  AOI22X1 U3095 ( .A(n8931), .B(recentABools_len_new_reg_385[28]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[28]), .D(n8657), .Y(n2344)
         );
  OAI21X1 U3096 ( .A(ap_CS_fsm[12]), .B(n10631), .C(n7919), .Y(n4313) );
  AOI22X1 U3097 ( .A(n8931), .B(recentABools_len_new_reg_385[27]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[27]), .D(n8657), .Y(n2346)
         );
  OAI21X1 U3098 ( .A(ap_CS_fsm[12]), .B(n10630), .C(n7702), .Y(n4314) );
  AOI22X1 U3099 ( .A(n8931), .B(recentABools_len_new_reg_385[26]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[26]), .D(n8657), .Y(n2348)
         );
  OAI21X1 U3101 ( .A(ap_CS_fsm[12]), .B(n10629), .C(n7501), .Y(n4315) );
  AOI22X1 U3102 ( .A(n8931), .B(recentABools_len_new_reg_385[25]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[25]), .D(n8657), .Y(n2350)
         );
  OAI21X1 U3104 ( .A(ap_CS_fsm[12]), .B(n10628), .C(n8164), .Y(n4316) );
  AOI22X1 U3105 ( .A(n8931), .B(recentABools_len_new_reg_385[24]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[24]), .D(n8657), .Y(n2352)
         );
  OAI21X1 U3106 ( .A(ap_CS_fsm[12]), .B(n10627), .C(n7322), .Y(n4317) );
  AOI22X1 U3107 ( .A(n8931), .B(recentABools_len_new_reg_385[23]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[23]), .D(n8657), .Y(n2354)
         );
  OAI21X1 U3108 ( .A(ap_CS_fsm[12]), .B(n10626), .C(n7158), .Y(n4318) );
  AOI22X1 U3109 ( .A(n8931), .B(recentABools_len_new_reg_385[22]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[22]), .D(n8657), .Y(n2356)
         );
  OAI21X1 U3111 ( .A(ap_CS_fsm[12]), .B(n10625), .C(n7009), .Y(n4319) );
  AOI22X1 U3112 ( .A(n8931), .B(recentABools_len_new_reg_385[21]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[21]), .D(n8657), .Y(n2358)
         );
  OAI21X1 U3114 ( .A(ap_CS_fsm[12]), .B(n10624), .C(n6868), .Y(n4320) );
  AOI22X1 U3115 ( .A(n8931), .B(recentABools_len_new_reg_385[20]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[20]), .D(n8657), .Y(n2360)
         );
  OAI21X1 U3117 ( .A(ap_CS_fsm[12]), .B(n10623), .C(n6740), .Y(n4321) );
  AOI22X1 U3118 ( .A(n8931), .B(recentABools_len_new_reg_385[19]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[19]), .D(n8657), .Y(n2362)
         );
  OAI21X1 U3120 ( .A(ap_CS_fsm[12]), .B(n10622), .C(n6622), .Y(n4322) );
  AOI22X1 U3121 ( .A(n8931), .B(recentABools_len_new_reg_385[18]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[18]), .D(n8657), .Y(n2364)
         );
  OAI21X1 U3122 ( .A(ap_CS_fsm[12]), .B(n10621), .C(n6510), .Y(n4323) );
  AOI22X1 U3123 ( .A(n8931), .B(recentABools_len_new_reg_385[17]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[17]), .D(n8657), .Y(n2366)
         );
  OAI21X1 U3124 ( .A(ap_CS_fsm[12]), .B(n10620), .C(n6403), .Y(n4324) );
  AOI22X1 U3125 ( .A(n8931), .B(recentABools_len_new_reg_385[16]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[16]), .D(n8657), .Y(n2368)
         );
  OAI21X1 U3126 ( .A(ap_CS_fsm[12]), .B(n10619), .C(n6297), .Y(n4325) );
  AOI22X1 U3127 ( .A(n8931), .B(recentABools_len_new_reg_385[15]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[15]), .D(n8657), .Y(n2370)
         );
  OAI21X1 U3128 ( .A(ap_CS_fsm[12]), .B(n10618), .C(n7918), .Y(n4326) );
  AOI22X1 U3129 ( .A(n8931), .B(recentABools_len_new_reg_385[14]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[14]), .D(n8657), .Y(n2372)
         );
  OAI21X1 U3130 ( .A(ap_CS_fsm[12]), .B(n10617), .C(n6204), .Y(n4327) );
  AOI22X1 U3131 ( .A(n8931), .B(recentABools_len_new_reg_385[13]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[13]), .D(n8657), .Y(n2374)
         );
  OAI21X1 U3132 ( .A(ap_CS_fsm[12]), .B(n10616), .C(n7701), .Y(n4328) );
  AOI22X1 U3133 ( .A(n8931), .B(recentABools_len_new_reg_385[12]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[12]), .D(n8657), .Y(n2376)
         );
  OAI21X1 U3134 ( .A(ap_CS_fsm[12]), .B(n10615), .C(n7499), .Y(n4329) );
  AOI22X1 U3135 ( .A(n8931), .B(recentABools_len_new_reg_385[11]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[11]), .D(n8657), .Y(n2378)
         );
  OAI21X1 U3136 ( .A(ap_CS_fsm[12]), .B(n10614), .C(n7156), .Y(n4330) );
  AOI22X1 U3137 ( .A(n8931), .B(recentABools_len_new_reg_385[10]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[10]), .D(n8657), .Y(n2380)
         );
  OAI21X1 U3139 ( .A(ap_CS_fsm[12]), .B(n10613), .C(n7320), .Y(n4331) );
  AOI22X1 U3140 ( .A(n8931), .B(recentABools_len_new_reg_385[9]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[9]), .D(n8657), .Y(n2382)
         );
  OAI21X1 U3142 ( .A(ap_CS_fsm[12]), .B(n10612), .C(n7007), .Y(n4332) );
  AOI22X1 U3143 ( .A(n8931), .B(recentABools_len_new_reg_385[8]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[8]), .D(n8657), .Y(n2384)
         );
  OAI21X1 U3145 ( .A(ap_CS_fsm[12]), .B(n10611), .C(n6866), .Y(n4333) );
  AOI22X1 U3146 ( .A(n8931), .B(recentABools_len_new_reg_385[7]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[7]), .D(n8657), .Y(n2386)
         );
  OAI21X1 U3147 ( .A(ap_CS_fsm[12]), .B(n10610), .C(n6738), .Y(n4334) );
  AOI22X1 U3148 ( .A(n8931), .B(recentABools_len_new_reg_385[6]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[6]), .D(n8657), .Y(n2388)
         );
  OAI21X1 U3149 ( .A(ap_CS_fsm[12]), .B(n10609), .C(n6620), .Y(n4335) );
  AOI22X1 U3150 ( .A(n8931), .B(recentABools_len_new_reg_385[5]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[5]), .D(n8657), .Y(n2390)
         );
  OAI21X1 U3151 ( .A(ap_CS_fsm[12]), .B(n10608), .C(n6508), .Y(n4336) );
  AOI22X1 U3152 ( .A(n8931), .B(recentABools_len_new_reg_385[4]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[4]), .D(n8657), .Y(n2392)
         );
  OAI21X1 U3153 ( .A(ap_CS_fsm[12]), .B(n10607), .C(n7917), .Y(n4337) );
  AOI22X1 U3154 ( .A(n8931), .B(recentABools_len_new_reg_385[3]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[3]), .D(n8657), .Y(n2394)
         );
  OAI21X1 U3155 ( .A(ap_CS_fsm[12]), .B(n10606), .C(n6401), .Y(n4338) );
  AOI22X1 U3156 ( .A(n8931), .B(recentABools_len_new_reg_385[2]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[2]), .D(n8657), .Y(n2396)
         );
  OAI21X1 U3158 ( .A(ap_CS_fsm[12]), .B(n10605), .C(n6295), .Y(n4339) );
  AOI22X1 U3159 ( .A(n8931), .B(recentABools_len_new_reg_385[1]), .C(n10574), 
        .D(n8657), .Y(n2398) );
  OAI21X1 U3161 ( .A(ap_CS_fsm[12]), .B(n10540), .C(n4805), .Y(n4340) );
  AOI22X1 U3162 ( .A(n8931), .B(recentABools_len_new_reg_385[0]), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[0]), .D(n8657), .Y(n2400)
         );
  OAI21X1 U3165 ( .A(n7095), .B(n2239), .C(n4804), .Y(n4341) );
  AOI22X1 U3166 ( .A(recentABools_len_new_reg_385[31]), .B(n8932), .C(
        CircularBuffer_len_write_assig_3_fu_1249_p2[31]), .D(n8890), .Y(n2402)
         );
  OAI21X1 U3171 ( .A(ap_CS_fsm[12]), .B(n10543), .C(n6200), .Y(n4342) );
  OAI21X1 U3173 ( .A(n8930), .B(n9382), .C(n6914), .Y(sum_1_phi_fu_379_p4[0])
         );
  OAI21X1 U3176 ( .A(ap_CS_fsm[12]), .B(n10544), .C(n6124), .Y(n4343) );
  OAI21X1 U3178 ( .A(n8930), .B(n9381), .C(n7212), .Y(sum_1_phi_fu_379_p4[1])
         );
  OAI21X1 U3181 ( .A(ap_CS_fsm[12]), .B(n10545), .C(n6615), .Y(n4344) );
  OAI21X1 U3183 ( .A(n8930), .B(n9379), .C(n7378), .Y(sum_1_phi_fu_379_p4[2])
         );
  OAI21X1 U3186 ( .A(ap_CS_fsm[12]), .B(n10546), .C(n6502), .Y(n4345) );
  OAI21X1 U3188 ( .A(n8930), .B(n9378), .C(n6659), .Y(sum_1_phi_fu_379_p4[3])
         );
  OAI21X1 U3191 ( .A(ap_CS_fsm[12]), .B(n10547), .C(n6732), .Y(n4346) );
  OAI21X1 U3193 ( .A(n8930), .B(n9375), .C(n8214), .Y(sum_1_phi_fu_379_p4[4])
         );
  OAI21X1 U3196 ( .A(ap_CS_fsm[12]), .B(n10548), .C(n6860), .Y(n4347) );
  OAI21X1 U3198 ( .A(n8930), .B(n9374), .C(n7758), .Y(sum_1_phi_fu_379_p4[5])
         );
  OAI21X1 U3201 ( .A(ap_CS_fsm[12]), .B(n10549), .C(n6999), .Y(n4348) );
  OAI21X1 U3203 ( .A(n8930), .B(n9373), .C(n7560), .Y(sum_1_phi_fu_379_p4[6])
         );
  OAI21X1 U3206 ( .A(ap_CS_fsm[12]), .B(n10550), .C(n6059), .Y(n4349) );
  OAI21X1 U3208 ( .A(n8930), .B(n9372), .C(n6152), .Y(sum_1_phi_fu_379_p4[7])
         );
  OAI21X1 U3211 ( .A(ap_CS_fsm[12]), .B(n10551), .C(n6202), .Y(n4350) );
  OAI21X1 U3213 ( .A(n8930), .B(n9369), .C(n6085), .Y(sum_1_phi_fu_379_p4[8])
         );
  OAI21X1 U3216 ( .A(ap_CS_fsm[12]), .B(n10552), .C(n6292), .Y(n4351) );
  OAI21X1 U3218 ( .A(n8930), .B(n9367), .C(n6916), .Y(sum_1_phi_fu_379_p4[9])
         );
  OAI21X1 U3221 ( .A(ap_CS_fsm[12]), .B(n10553), .C(n6504), .Y(n4352) );
  OAI21X1 U3223 ( .A(n8930), .B(n9365), .C(n6783), .Y(sum_1_phi_fu_379_p4[10])
         );
  OAI21X1 U3226 ( .A(ap_CS_fsm[12]), .B(n10554), .C(n6397), .Y(n4353) );
  OAI21X1 U3228 ( .A(n8930), .B(n9364), .C(n5053), .Y(sum_1_phi_fu_379_p4[11])
         );
  OAI21X1 U3231 ( .A(ap_CS_fsm[12]), .B(n10555), .C(n6616), .Y(n4354) );
  OAI21X1 U3233 ( .A(n8930), .B(n9360), .C(n6439), .Y(sum_1_phi_fu_379_p4[12])
         );
  OAI21X1 U3236 ( .A(ap_CS_fsm[12]), .B(n10556), .C(n6733), .Y(n4355) );
  OAI21X1 U3238 ( .A(n8930), .B(n9359), .C(n6550), .Y(sum_1_phi_fu_379_p4[13])
         );
  OAI21X1 U3241 ( .A(ap_CS_fsm[12]), .B(n10557), .C(n6861), .Y(n4356) );
  OAI21X1 U3243 ( .A(n8930), .B(n9358), .C(n7063), .Y(sum_1_phi_fu_379_p4[14])
         );
  OAI21X1 U3246 ( .A(ap_CS_fsm[12]), .B(n10558), .C(n7150), .Y(n4357) );
  OAI21X1 U3248 ( .A(n8930), .B(n9357), .C(n6437), .Y(sum_1_phi_fu_379_p4[15])
         );
  OAI21X1 U3251 ( .A(ap_CS_fsm[12]), .B(n10559), .C(n7001), .Y(n4358) );
  OAI21X1 U3253 ( .A(n8930), .B(n9351), .C(n6661), .Y(sum_1_phi_fu_379_p4[16])
         );
  OAI21X1 U3256 ( .A(ap_CS_fsm[12]), .B(n10560), .C(n7314), .Y(n4359) );
  OAI21X1 U3258 ( .A(n8930), .B(n9350), .C(n8215), .Y(sum_1_phi_fu_379_p4[17])
         );
  OAI21X1 U3261 ( .A(ap_CS_fsm[12]), .B(n10561), .C(n7494), .Y(n4360) );
  OAI21X1 U3263 ( .A(n8930), .B(n9349), .C(n7760), .Y(sum_1_phi_fu_379_p4[18])
         );
  OAI21X1 U3266 ( .A(ap_CS_fsm[12]), .B(n10562), .C(n7697), .Y(n4361) );
  OAI21X1 U3268 ( .A(n8930), .B(n9348), .C(n5052), .Y(sum_1_phi_fu_379_p4[19])
         );
  OAI21X1 U3271 ( .A(ap_CS_fsm[12]), .B(n10563), .C(n7913), .Y(n4362) );
  OAI21X1 U3273 ( .A(n8930), .B(n9344), .C(n6781), .Y(sum_1_phi_fu_379_p4[20])
         );
  OAI21X1 U3276 ( .A(ap_CS_fsm[12]), .B(n10564), .C(n8162), .Y(n4363) );
  OAI21X1 U3278 ( .A(n8930), .B(n9343), .C(n7562), .Y(sum_1_phi_fu_379_p4[21])
         );
  OAI21X1 U3281 ( .A(ap_CS_fsm[12]), .B(n10565), .C(n6399), .Y(n4364) );
  OAI21X1 U3283 ( .A(n8930), .B(n9342), .C(n7978), .Y(sum_1_phi_fu_379_p4[22])
         );
  OAI21X1 U3286 ( .A(ap_CS_fsm[12]), .B(n10566), .C(n6506), .Y(n4365) );
  OAI21X1 U3288 ( .A(n8930), .B(n9341), .C(n6913), .Y(sum_1_phi_fu_379_p4[23])
         );
  OAI21X1 U3291 ( .A(ap_CS_fsm[12]), .B(n10567), .C(n6618), .Y(n4366) );
  OAI21X1 U3293 ( .A(n8930), .B(n9336), .C(n6330), .Y(sum_1_phi_fu_379_p4[24])
         );
  OAI21X1 U3296 ( .A(ap_CS_fsm[12]), .B(n10568), .C(n6735), .Y(n4367) );
  OAI21X1 U3298 ( .A(n8930), .B(n9335), .C(n7377), .Y(sum_1_phi_fu_379_p4[25])
         );
  OAI21X1 U3301 ( .A(ap_CS_fsm[12]), .B(n10569), .C(n6863), .Y(n4368) );
  OAI21X1 U3303 ( .A(n8930), .B(n9334), .C(n7219), .Y(sum_1_phi_fu_379_p4[26])
         );
  OAI21X1 U3306 ( .A(ap_CS_fsm[12]), .B(n10570), .C(n7003), .Y(n4369) );
  OAI21X1 U3308 ( .A(n8930), .B(n9333), .C(n6237), .Y(sum_1_phi_fu_379_p4[27])
         );
  OAI21X1 U3311 ( .A(ap_CS_fsm[12]), .B(n10571), .C(n7151), .Y(n4370) );
  OAI21X1 U3313 ( .A(n8930), .B(n9329), .C(n6327), .Y(sum_1_phi_fu_379_p4[28])
         );
  OAI21X1 U3316 ( .A(ap_CS_fsm[12]), .B(n10572), .C(n7316), .Y(n4371) );
  OAI21X1 U3318 ( .A(n8930), .B(n9328), .C(n7976), .Y(sum_1_phi_fu_379_p4[29])
         );
  OAI21X1 U3321 ( .A(ap_CS_fsm[12]), .B(n10811), .C(n7520), .Y(n4372) );
  OAI21X1 U3323 ( .A(n8930), .B(n9327), .C(n7058), .Y(sum_1_phi_fu_379_p4[30])
         );
  OAI21X1 U3326 ( .A(ap_CS_fsm[12]), .B(n9384), .C(n6255), .Y(n4373) );
  OAI21X1 U3328 ( .A(n8930), .B(n9326), .C(n6548), .Y(sum_1_phi_fu_379_p4[31])
         );
  OAI21X1 U3332 ( .A(n10532), .B(n2533), .C(n7695), .Y(n4374) );
  OAI21X1 U3335 ( .A(n10528), .B(n2533), .C(n8159), .Y(n4375) );
  OAI21X1 U3338 ( .A(n10526), .B(n2533), .C(n7492), .Y(n4376) );
  OAI21X1 U3341 ( .A(n10524), .B(n2533), .C(n7312), .Y(n4377) );
  OAI21X1 U3344 ( .A(n10522), .B(n2533), .C(n7910), .Y(n4378) );
  OAI21X1 U3347 ( .A(n10518), .B(n2533), .C(n7147), .Y(n4379) );
  OAI21X1 U3350 ( .A(n10516), .B(n2533), .C(n6998), .Y(n4380) );
  OAI21X1 U3353 ( .A(n10513), .B(n2533), .C(n6858), .Y(n4381) );
  OAI21X1 U3356 ( .A(n10511), .B(n2533), .C(n6730), .Y(n4382) );
  OAI21X1 U3359 ( .A(n10507), .B(n2533), .C(n6613), .Y(n4383) );
  OAI21X1 U3362 ( .A(n10505), .B(n2533), .C(n6501), .Y(n4384) );
  OAI21X1 U3365 ( .A(n10502), .B(n2533), .C(n6394), .Y(n4385) );
  OAI21X1 U3368 ( .A(n10500), .B(n2533), .C(n8156), .Y(n4386) );
  OAI21X1 U3371 ( .A(n10496), .B(n2533), .C(n7907), .Y(n4387) );
  OAI21X1 U3374 ( .A(n10494), .B(n2533), .C(n7308), .Y(n4388) );
  OAI21X1 U3377 ( .A(n10492), .B(n2533), .C(n7144), .Y(n4389) );
  OAI21X1 U3380 ( .A(n10490), .B(n2533), .C(n7691), .Y(n4390) );
  OAI21X1 U3383 ( .A(n10486), .B(n2533), .C(n7488), .Y(n4391) );
  OAI21X1 U3386 ( .A(n10484), .B(n2533), .C(n6995), .Y(n4392) );
  OAI21X1 U3389 ( .A(n10481), .B(n2533), .C(n6855), .Y(n4393) );
  OAI21X1 U3392 ( .A(n10479), .B(n2533), .C(n6727), .Y(n4394) );
  OAI21X1 U3395 ( .A(n10475), .B(n2533), .C(n6498), .Y(n4395) );
  OAI21X1 U3398 ( .A(n10473), .B(n2533), .C(n6609), .Y(n4396) );
  OAI21X1 U3401 ( .A(n10469), .B(n2533), .C(n6391), .Y(n4397) );
  OAI21X1 U3404 ( .A(n10467), .B(n2533), .C(n8154), .Y(n4398) );
  OAI21X1 U3407 ( .A(n10464), .B(n2533), .C(n7905), .Y(n4399) );
  OAI21X1 U3410 ( .A(n10462), .B(n2533), .C(n7487), .Y(n4400) );
  OAI21X1 U3413 ( .A(n10460), .B(n2533), .C(n7306), .Y(n4401) );
  OAI21X1 U3416 ( .A(n10458), .B(n2533), .C(n7689), .Y(n4402) );
  OAI21X1 U3419 ( .A(n10455), .B(n2533), .C(n7142), .Y(n4403) );
  OAI21X1 U3422 ( .A(n10453), .B(n2533), .C(n6993), .Y(n4404) );
  OAI21X1 U3425 ( .A(n10450), .B(n2533), .C(n6853), .Y(n4405) );
  OAI21X1 U3428 ( .A(\last_sample_is_V_V[0] ), .B(n9649), .C(ap_CS_fsm[7]), 
        .Y(n2533) );
  OAI21X1 U3431 ( .A(ap_CS_fsm[7]), .B(n10239), .C(n8378), .Y(n4406) );
  OAI21X1 U3433 ( .A(ap_CS_fsm[7]), .B(n10240), .C(n8378), .Y(n4407) );
  OAI21X1 U3436 ( .A(n9012), .B(n10241), .C(n7892), .Y(n4408) );
  OAI21X1 U3438 ( .A(n8929), .B(n10173), .C(n8209), .Y(sum_phi_fu_311_p4[31])
         );
  OAI21X1 U3441 ( .A(n9012), .B(n10238), .C(n7294), .Y(n4409) );
  OAI21X1 U3443 ( .A(n8929), .B(n10174), .C(n7553), .Y(sum_phi_fu_311_p4[30])
         );
  OAI21X1 U3446 ( .A(ap_CS_fsm[7]), .B(n10237), .C(n8144), .Y(n4410) );
  OAI21X1 U3448 ( .A(n8929), .B(n10175), .C(n7975), .Y(sum_phi_fu_311_p4[29])
         );
  OAI21X1 U3451 ( .A(n9012), .B(n10236), .C(n7472), .Y(n4411) );
  OAI21X1 U3453 ( .A(n8929), .B(n10176), .C(n6658), .Y(sum_phi_fu_311_p4[28])
         );
  OAI21X1 U3456 ( .A(n9012), .B(n10235), .C(n7129), .Y(n4412) );
  OAI21X1 U3458 ( .A(n8929), .B(n10177), .C(n7750), .Y(sum_phi_fu_311_p4[27])
         );
  OAI21X1 U3461 ( .A(ap_CS_fsm[7]), .B(n10234), .C(n8143), .Y(n4413) );
  OAI21X1 U3463 ( .A(n8929), .B(n10178), .C(n6786), .Y(sum_phi_fu_311_p4[26])
         );
  OAI21X1 U3466 ( .A(n9012), .B(n10233), .C(n6979), .Y(n4414) );
  OAI21X1 U3468 ( .A(n8929), .B(n10179), .C(n6921), .Y(sum_phi_fu_311_p4[25])
         );
  OAI21X1 U3471 ( .A(n9012), .B(n10232), .C(n6840), .Y(n4415) );
  OAI21X1 U3473 ( .A(n8929), .B(n10180), .C(n6438), .Y(sum_phi_fu_311_p4[24])
         );
  OAI21X1 U3476 ( .A(ap_CS_fsm[7]), .B(n10231), .C(n6712), .Y(n4416) );
  OAI21X1 U3478 ( .A(n8929), .B(n10181), .C(n6151), .Y(sum_phi_fu_311_p4[23])
         );
  OAI21X1 U3481 ( .A(ap_CS_fsm[7]), .B(n10230), .C(n6595), .Y(n4417) );
  OAI21X1 U3483 ( .A(n8929), .B(n10182), .C(n7064), .Y(sum_phi_fu_311_p4[22])
         );
  OAI21X1 U3486 ( .A(n9012), .B(n10229), .C(n6484), .Y(n4418) );
  OAI21X1 U3488 ( .A(n8929), .B(n10183), .C(n7376), .Y(sum_phi_fu_311_p4[21])
         );
  OAI21X1 U3491 ( .A(n9012), .B(n10228), .C(n6377), .Y(n4419) );
  OAI21X1 U3493 ( .A(n8929), .B(n10184), .C(n6329), .Y(sum_phi_fu_311_p4[20])
         );
  OAI21X1 U3496 ( .A(n9012), .B(n10227), .C(n6275), .Y(n4420) );
  OAI21X1 U3498 ( .A(n8929), .B(n10185), .C(n5051), .Y(sum_phi_fu_311_p4[19])
         );
  OAI21X1 U3501 ( .A(n9012), .B(n10226), .C(n6186), .Y(n4421) );
  OAI21X1 U3503 ( .A(n8929), .B(n10186), .C(n7977), .Y(sum_phi_fu_311_p4[18])
         );
  OAI21X1 U3506 ( .A(n9012), .B(n10225), .C(n6112), .Y(n4422) );
  OAI21X1 U3508 ( .A(n8929), .B(n10187), .C(n7220), .Y(sum_phi_fu_311_p4[17])
         );
  OAI21X1 U3511 ( .A(n9012), .B(n10224), .C(n7890), .Y(n4423) );
  OAI21X1 U3513 ( .A(n8929), .B(n10188), .C(n7379), .Y(sum_phi_fu_311_p4[16])
         );
  OAI21X1 U3516 ( .A(n9012), .B(n10223), .C(n7675), .Y(n4424) );
  OAI21X1 U3518 ( .A(n8929), .B(n10189), .C(n6236), .Y(sum_phi_fu_311_p4[15])
         );
  OAI21X1 U3521 ( .A(n9012), .B(n10222), .C(n7292), .Y(n4425) );
  OAI21X1 U3523 ( .A(n8929), .B(n10190), .C(n6915), .Y(sum_phi_fu_311_p4[14])
         );
  OAI21X1 U3526 ( .A(n9012), .B(n10221), .C(n7470), .Y(n4426) );
  OAI21X1 U3528 ( .A(n8929), .B(n10191), .C(n6779), .Y(sum_phi_fu_311_p4[13])
         );
  OAI21X1 U3531 ( .A(ap_CS_fsm[7]), .B(n10220), .C(n7126), .Y(n4427) );
  OAI21X1 U3533 ( .A(n8929), .B(n10192), .C(n6549), .Y(sum_phi_fu_311_p4[12])
         );
  OAI21X1 U3536 ( .A(n9012), .B(n10219), .C(n6977), .Y(n4428) );
  OAI21X1 U3538 ( .A(n8929), .B(n10193), .C(n6436), .Y(sum_phi_fu_311_p4[11])
         );
  OAI21X1 U3541 ( .A(n9012), .B(n10218), .C(n6837), .Y(n4429) );
  OAI21X1 U3543 ( .A(n8929), .B(n10194), .C(n7057), .Y(sum_phi_fu_311_p4[10])
         );
  OAI21X1 U3546 ( .A(n9012), .B(n10217), .C(n6594), .Y(n4430) );
  OAI21X1 U3548 ( .A(n8929), .B(n10195), .C(n7561), .Y(sum_phi_fu_311_p4[9])
         );
  OAI21X1 U3551 ( .A(ap_CS_fsm[7]), .B(n10216), .C(n6710), .Y(n4431) );
  OAI21X1 U3553 ( .A(n8929), .B(n10196), .C(n7968), .Y(sum_phi_fu_311_p4[8])
         );
  OAI21X1 U3556 ( .A(ap_CS_fsm[7]), .B(n10215), .C(n6482), .Y(n4432) );
  OAI21X1 U3558 ( .A(n8929), .B(n10197), .C(n6084), .Y(sum_phi_fu_311_p4[7])
         );
  OAI21X1 U3561 ( .A(ap_CS_fsm[7]), .B(n10214), .C(n6374), .Y(n4433) );
  OAI21X1 U3563 ( .A(n8929), .B(n10198), .C(n7759), .Y(sum_phi_fu_311_p4[6])
         );
  OAI21X1 U3566 ( .A(ap_CS_fsm[7]), .B(n10213), .C(n6273), .Y(n4434) );
  OAI21X1 U3568 ( .A(n8929), .B(n10199), .C(n8213), .Y(sum_phi_fu_311_p4[5])
         );
  OAI21X1 U3571 ( .A(n9012), .B(n10212), .C(n6184), .Y(n4435) );
  OAI21X1 U3573 ( .A(n8929), .B(n10200), .C(n6660), .Y(sum_phi_fu_311_p4[4])
         );
  OAI21X1 U3576 ( .A(ap_CS_fsm[7]), .B(n10211), .C(n6110), .Y(n4436) );
  OAI21X1 U3578 ( .A(n8929), .B(n10201), .C(n7211), .Y(sum_phi_fu_311_p4[3])
         );
  OAI21X1 U3581 ( .A(ap_CS_fsm[7]), .B(n10210), .C(n6049), .Y(n4437) );
  OAI21X1 U3583 ( .A(n8929), .B(n10202), .C(n6328), .Y(sum_phi_fu_311_p4[2])
         );
  OAI21X1 U3586 ( .A(ap_CS_fsm[7]), .B(n10209), .C(n7889), .Y(n4438) );
  OAI21X1 U3588 ( .A(n8929), .B(n10203), .C(n6547), .Y(sum_phi_fu_311_p4[1])
         );
  OAI21X1 U3591 ( .A(n9012), .B(n10208), .C(n8142), .Y(n4439) );
  OAI21X1 U3593 ( .A(n8929), .B(n10204), .C(n6235), .Y(sum_phi_fu_311_p4[0])
         );
  OAI21X1 U3596 ( .A(n4688), .B(n8927), .C(n7891), .Y(n4440) );
  AOI22X1 U3597 ( .A(n8925), .B(sum_reg_308[31]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[31]), .Y(n2700) );
  OAI21X1 U3599 ( .A(n8459), .B(n8927), .C(n7677), .Y(n4441) );
  AOI22X1 U3600 ( .A(n8925), .B(sum_reg_308[30]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[30]), .Y(n2703) );
  OAI21X1 U3602 ( .A(n8460), .B(n8927), .C(n7473), .Y(n4442) );
  AOI22X1 U3603 ( .A(n8925), .B(sum_reg_308[29]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[29]), .Y(n2704) );
  OAI21X1 U3605 ( .A(n8461), .B(n8927), .C(n7293), .Y(n4443) );
  AOI22X1 U3606 ( .A(n8925), .B(sum_reg_308[28]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[28]), .Y(n2705) );
  OAI21X1 U3608 ( .A(n8462), .B(n8927), .C(n7128), .Y(n4444) );
  AOI22X1 U3609 ( .A(n8925), .B(sum_reg_308[27]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[27]), .Y(n2706) );
  OAI21X1 U3611 ( .A(n8463), .B(n8927), .C(n6980), .Y(n4445) );
  AOI22X1 U3612 ( .A(n8925), .B(sum_reg_308[26]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[26]), .Y(n2707) );
  OAI21X1 U3614 ( .A(n8464), .B(n2699), .C(n6713), .Y(n4446) );
  AOI22X1 U3615 ( .A(n8925), .B(sum_reg_308[25]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[25]), .Y(n2708) );
  OAI21X1 U3617 ( .A(n8465), .B(n8927), .C(n6839), .Y(n4447) );
  AOI22X1 U3618 ( .A(n8925), .B(sum_reg_308[24]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[24]), .Y(n2709) );
  OAI21X1 U3620 ( .A(n8466), .B(n2699), .C(n6596), .Y(n4448) );
  AOI22X1 U3621 ( .A(n8925), .B(sum_reg_308[23]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[23]), .Y(n2710) );
  OAI21X1 U3623 ( .A(n8467), .B(n8927), .C(n6485), .Y(n4449) );
  AOI22X1 U3624 ( .A(n8925), .B(sum_reg_308[22]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[22]), .Y(n2711) );
  OAI21X1 U3626 ( .A(n8468), .B(n2699), .C(n6276), .Y(n4450) );
  AOI22X1 U3627 ( .A(n8925), .B(sum_reg_308[21]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[21]), .Y(n2712) );
  OAI21X1 U3629 ( .A(n8469), .B(n8927), .C(n6376), .Y(n4451) );
  AOI22X1 U3630 ( .A(n8925), .B(sum_reg_308[20]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[20]), .Y(n2713) );
  OAI21X1 U3632 ( .A(n8470), .B(n8927), .C(n6187), .Y(n4452) );
  AOI22X1 U3633 ( .A(n8925), .B(sum_reg_308[19]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[19]), .Y(n2714) );
  OAI21X1 U3635 ( .A(n8471), .B(n2699), .C(n6113), .Y(n4453) );
  AOI22X1 U3636 ( .A(n2701), .B(sum_reg_308[18]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[18]), .Y(n2715) );
  OAI21X1 U3638 ( .A(n8472), .B(n2699), .C(n7676), .Y(n4454) );
  AOI22X1 U3639 ( .A(n8925), .B(sum_reg_308[17]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[17]), .Y(n2716) );
  OAI21X1 U3641 ( .A(n8473), .B(n8927), .C(n7471), .Y(n4455) );
  AOI22X1 U3642 ( .A(n2701), .B(sum_reg_308[16]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[16]), .Y(n2717) );
  OAI21X1 U3644 ( .A(n8474), .B(n8927), .C(n7127), .Y(n4456) );
  AOI22X1 U3645 ( .A(n8925), .B(sum_reg_308[15]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[15]), .Y(n2718) );
  OAI21X1 U3647 ( .A(n8475), .B(n2699), .C(n7291), .Y(n4457) );
  AOI22X1 U3648 ( .A(n2701), .B(sum_reg_308[14]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[14]), .Y(n2719) );
  OAI21X1 U3650 ( .A(n8476), .B(n8927), .C(n6978), .Y(n4458) );
  AOI22X1 U3651 ( .A(n8925), .B(sum_reg_308[13]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[13]), .Y(n2720) );
  OAI21X1 U3653 ( .A(n8477), .B(n8927), .C(n6838), .Y(n4459) );
  AOI22X1 U3654 ( .A(n2701), .B(sum_reg_308[12]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[12]), .Y(n2721) );
  OAI21X1 U3656 ( .A(n8478), .B(n8927), .C(n6711), .Y(n4460) );
  AOI22X1 U3657 ( .A(n8925), .B(sum_reg_308[11]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[11]), .Y(n2722) );
  OAI21X1 U3659 ( .A(n8479), .B(n2699), .C(n6483), .Y(n4461) );
  AOI22X1 U3660 ( .A(n2701), .B(sum_reg_308[10]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[10]), .Y(n2723) );
  OAI21X1 U3662 ( .A(n8480), .B(n8927), .C(n6593), .Y(n4462) );
  AOI22X1 U3663 ( .A(n8925), .B(sum_reg_308[9]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[9]), .Y(n2724) );
  OAI21X1 U3665 ( .A(n8481), .B(n8927), .C(n6375), .Y(n4463) );
  AOI22X1 U3666 ( .A(n2701), .B(sum_reg_308[8]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[8]), .Y(n2725) );
  OAI21X1 U3668 ( .A(n8482), .B(n2699), .C(n6274), .Y(n4464) );
  AOI22X1 U3669 ( .A(n8925), .B(sum_reg_308[7]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[7]), .Y(n2726) );
  OAI21X1 U3671 ( .A(n8483), .B(n2699), .C(n6185), .Y(n4465) );
  AOI22X1 U3672 ( .A(n2701), .B(sum_reg_308[6]), .C(n2864), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[6]), .Y(n2727) );
  OAI21X1 U3674 ( .A(n8484), .B(n8927), .C(n6111), .Y(n4466) );
  AOI22X1 U3675 ( .A(n2701), .B(sum_reg_308[5]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[5]), .Y(n2728) );
  OAI21X1 U3677 ( .A(n8485), .B(n8927), .C(n7674), .Y(n4467) );
  AOI22X1 U3678 ( .A(n8925), .B(sum_reg_308[4]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[4]), .Y(n2729) );
  OAI21X1 U3680 ( .A(n8486), .B(n2699), .C(n7469), .Y(n4468) );
  AOI22X1 U3681 ( .A(n8925), .B(sum_reg_308[3]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[3]), .Y(n2730) );
  OAI21X1 U3683 ( .A(n8487), .B(n8927), .C(n7290), .Y(n4469) );
  AOI22X1 U3684 ( .A(n2701), .B(sum_reg_308[2]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[2]), .Y(n2731) );
  OAI21X1 U3686 ( .A(n8488), .B(n2699), .C(n7125), .Y(n4470) );
  AOI22X1 U3687 ( .A(n2701), .B(sum_reg_308[1]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[1]), .Y(n2732) );
  OAI21X1 U3689 ( .A(n8663), .B(n8927), .C(n6976), .Y(n4471) );
  AOI22X1 U3690 ( .A(n8925), .B(sum_reg_308[0]), .C(n8893), .D(
        CircularBuffer_sum_write_assig_1_fu_917_p2[0]), .Y(n2733) );
  OAI21X1 U3692 ( .A(n7259), .B(n2699), .C(n6177), .Y(n4472) );
  AOI22X1 U3693 ( .A(recentVBools_len_new_reg_317[30]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[30]), .D(n8893), .Y(n2735)
         );
  OAI21X1 U3694 ( .A(n6165), .B(n8927), .C(n4803), .Y(n4473) );
  AOI22X1 U3695 ( .A(recentVBools_len_new_reg_317[29]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[29]), .D(n8893), .Y(n2737)
         );
  OAI21X1 U3696 ( .A(n6687), .B(n8927), .C(n4802), .Y(n4474) );
  AOI22X1 U3697 ( .A(recentVBools_len_new_reg_317[28]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[28]), .D(n8893), .Y(n2739)
         );
  OAI21X1 U3698 ( .A(n7645), .B(n2699), .C(n6832), .Y(n4475) );
  AOI22X1 U3699 ( .A(recentVBools_len_new_reg_317[27]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[27]), .D(n8893), .Y(n2741)
         );
  OAI21X1 U3700 ( .A(n6812), .B(n8927), .C(n6478), .Y(n4476) );
  AOI22X1 U3701 ( .A(recentVBools_len_new_reg_317[26]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[26]), .D(n8893), .Y(n2743)
         );
  OAI21X1 U3702 ( .A(n6947), .B(n8927), .C(n6704), .Y(n4477) );
  AOI22X1 U3703 ( .A(recentVBools_len_new_reg_317[25]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[25]), .D(n8893), .Y(n2745)
         );
  OAI21X1 U3704 ( .A(n6572), .B(n2699), .C(n6370), .Y(n4478) );
  AOI22X1 U3705 ( .A(recentVBools_len_new_reg_317[24]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[24]), .D(n8893), .Y(n2747)
         );
  OAI21X1 U3706 ( .A(n8400), .B(n8927), .C(n6588), .Y(n4479) );
  AOI22X1 U3707 ( .A(recentVBools_len_new_reg_317[23]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[23]), .D(n8893), .Y(n2749)
         );
  OAI21X1 U3708 ( .A(n7099), .B(n8927), .C(n4801), .Y(n4480) );
  AOI22X1 U3709 ( .A(recentVBools_len_new_reg_317[22]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[22]), .D(n2864), .Y(n2751)
         );
  OAI21X1 U3710 ( .A(n7264), .B(n8927), .C(n4800), .Y(n4481) );
  AOI22X1 U3711 ( .A(recentVBools_len_new_reg_317[21]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[21]), .D(n2864), .Y(n2753)
         );
  OAI21X1 U3712 ( .A(n6459), .B(n8927), .C(n4799), .Y(n4482) );
  AOI22X1 U3713 ( .A(recentVBools_len_new_reg_317[20]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[20]), .D(n2864), .Y(n2755)
         );
  OAI21X1 U3714 ( .A(n7863), .B(n8927), .C(n7463), .Y(n4483) );
  AOI22X1 U3715 ( .A(recentVBools_len_new_reg_317[19]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[19]), .D(n2864), .Y(n2757)
         );
  OAI21X1 U3716 ( .A(n7442), .B(n8927), .C(n7121), .Y(n4484) );
  AOI22X1 U3717 ( .A(recentVBools_len_new_reg_317[18]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[18]), .D(n2864), .Y(n2759)
         );
  OAI21X1 U3718 ( .A(n6350), .B(n8927), .C(n4798), .Y(n4485) );
  AOI22X1 U3719 ( .A(recentVBools_len_new_reg_317[17]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[17]), .D(n2864), .Y(n2761)
         );
  OAI21X1 U3720 ( .A(n6253), .B(n8927), .C(n4797), .Y(n4486) );
  AOI22X1 U3721 ( .A(recentVBools_len_new_reg_317[16]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[16]), .D(n2864), .Y(n2763)
         );
  OAI21X1 U3722 ( .A(n8113), .B(n8927), .C(n7284), .Y(n4487) );
  AOI22X1 U3723 ( .A(recentVBools_len_new_reg_317[15]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[15]), .D(n2864), .Y(n2765)
         );
  OAI21X1 U3724 ( .A(n8102), .B(n8927), .C(n6970), .Y(n4488) );
  AOI22X1 U3725 ( .A(recentVBools_len_new_reg_317[14]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[14]), .D(n2864), .Y(n2767)
         );
  OAI21X1 U3726 ( .A(n7641), .B(n8927), .C(n6831), .Y(n4489) );
  AOI22X1 U3727 ( .A(recentVBools_len_new_reg_317[13]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[13]), .D(n2864), .Y(n2769)
         );
  OAI21X1 U3728 ( .A(n7438), .B(n2699), .C(n6269), .Y(n4490) );
  AOI22X1 U3729 ( .A(recentVBools_len_new_reg_317[12]), .B(n8925), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[12]), .D(n2864), .Y(n2771)
         );
  OAI21X1 U3730 ( .A(n8398), .B(n8927), .C(n6703), .Y(n4491) );
  AOI22X1 U3731 ( .A(recentVBools_len_new_reg_317[11]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[11]), .D(n2864), .Y(n2773)
         );
  OAI21X1 U3732 ( .A(n7859), .B(n8927), .C(n6587), .Y(n4492) );
  AOI22X1 U3733 ( .A(recentVBools_len_new_reg_317[10]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[10]), .D(n8893), .Y(n2775)
         );
  OAI21X1 U3734 ( .A(n7861), .B(n2699), .C(n7119), .Y(n4493) );
  AOI22X1 U3735 ( .A(recentVBools_len_new_reg_317[9]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[9]), .D(n2864), .Y(n2777)
         );
  OAI21X1 U3736 ( .A(n8406), .B(n2699), .C(n7462), .Y(n4494) );
  AOI22X1 U3737 ( .A(recentVBools_len_new_reg_317[8]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[8]), .D(n8893), .Y(n2779)
         );
  OAI21X1 U3738 ( .A(n8111), .B(n2699), .C(n7283), .Y(n4495) );
  AOI22X1 U3739 ( .A(recentVBools_len_new_reg_317[7]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[7]), .D(n2864), .Y(n2781)
         );
  OAI21X1 U3740 ( .A(n7643), .B(n2699), .C(n6968), .Y(n4496) );
  AOI22X1 U3741 ( .A(recentVBools_len_new_reg_317[6]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[6]), .D(n8893), .Y(n2783)
         );
  OAI21X1 U3742 ( .A(n7440), .B(n2699), .C(n6829), .Y(n4497) );
  AOI22X1 U3743 ( .A(recentVBools_len_new_reg_317[5]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[5]), .D(n2864), .Y(n2785)
         );
  OAI21X1 U3744 ( .A(n10071), .B(n2699), .C(n6701), .Y(n4498) );
  AOI22X1 U3745 ( .A(recentVBools_len_new_reg_317[4]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[4]), .D(n8893), .Y(n2787)
         );
  OAI21X1 U3747 ( .A(n10072), .B(n2699), .C(n6475), .Y(n4499) );
  AOI22X1 U3748 ( .A(recentVBools_len_new_reg_317[3]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[3]), .D(n2864), .Y(n2789)
         );
  OAI21X1 U3750 ( .A(n10073), .B(n8927), .C(n6367), .Y(n4500) );
  AOI22X1 U3751 ( .A(recentVBools_len_new_reg_317[2]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[2]), .D(n8893), .Y(n2791)
         );
  OAI21X1 U3753 ( .A(n10074), .B(n2699), .C(n6267), .Y(n4501) );
  AOI22X1 U3754 ( .A(recentVBools_len_new_reg_317[1]), .B(n2701), .C(n10079), 
        .D(n2864), .Y(n2793) );
  OAI21X1 U3756 ( .A(n8391), .B(n8927), .C(n7671), .Y(n4502) );
  AOI22X1 U3757 ( .A(recentVBools_len_new_reg_317[0]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[0]), .D(n8893), .Y(n2795)
         );
  OAI21X1 U3758 ( .A(n9012), .B(n10172), .C(n7670), .Y(n4503) );
  AOI22X1 U3759 ( .A(recentVBools_len_new_reg_317[31]), .B(n8924), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[31]), .D(n8656), .Y(n2797)
         );
  OAI21X1 U3760 ( .A(ap_CS_fsm[7]), .B(n10078), .C(n6364), .Y(n4504) );
  AOI22X1 U3761 ( .A(n8924), .B(recentVBools_len_new_reg_317[30]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[30]), .D(n8656), .Y(n2801)
         );
  OAI21X1 U3762 ( .A(ap_CS_fsm[7]), .B(n10138), .C(n8137), .Y(n4505) );
  AOI22X1 U3763 ( .A(n8924), .B(recentVBools_len_new_reg_317[29]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[29]), .D(n8656), .Y(n2803)
         );
  OAI21X1 U3764 ( .A(ap_CS_fsm[7]), .B(n10137), .C(n7885), .Y(n4506) );
  AOI22X1 U3765 ( .A(n8924), .B(recentVBools_len_new_reg_317[28]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[28]), .D(n8656), .Y(n2805)
         );
  OAI21X1 U3766 ( .A(n9012), .B(n10136), .C(n6705), .Y(n4507) );
  AOI22X1 U3767 ( .A(n8924), .B(recentVBools_len_new_reg_317[27]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[27]), .D(n8656), .Y(n2807)
         );
  OAI21X1 U3768 ( .A(ap_CS_fsm[7]), .B(n10135), .C(n6589), .Y(n4508) );
  AOI22X1 U3769 ( .A(n8924), .B(recentVBools_len_new_reg_317[26]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[26]), .D(n8656), .Y(n2809)
         );
  OAI21X1 U3771 ( .A(ap_CS_fsm[7]), .B(n10134), .C(n6477), .Y(n4509) );
  AOI22X1 U3772 ( .A(n8924), .B(recentVBools_len_new_reg_317[25]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[25]), .D(n8656), .Y(n2811)
         );
  OAI21X1 U3774 ( .A(n9012), .B(n10133), .C(n8136), .Y(n4510) );
  AOI22X1 U3775 ( .A(n8924), .B(recentVBools_len_new_reg_317[24]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[24]), .D(n8656), .Y(n2813)
         );
  OAI21X1 U3776 ( .A(n9012), .B(n10132), .C(n7668), .Y(n4511) );
  AOI22X1 U3777 ( .A(n8924), .B(recentVBools_len_new_reg_317[23]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[23]), .D(n8656), .Y(n2815)
         );
  OAI21X1 U3778 ( .A(n9012), .B(n10131), .C(n7285), .Y(n4512) );
  AOI22X1 U3779 ( .A(n8924), .B(recentVBools_len_new_reg_317[22]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[22]), .D(n8656), .Y(n2817)
         );
  OAI21X1 U3781 ( .A(n9012), .B(n10130), .C(n7122), .Y(n4513) );
  AOI22X1 U3782 ( .A(n8924), .B(recentVBools_len_new_reg_317[21]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[21]), .D(n8656), .Y(n2819)
         );
  OAI21X1 U3784 ( .A(n9012), .B(n10129), .C(n7464), .Y(n4514) );
  AOI22X1 U3785 ( .A(n8924), .B(recentVBools_len_new_reg_317[20]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[20]), .D(n8656), .Y(n2821)
         );
  OAI21X1 U3787 ( .A(n9012), .B(n10128), .C(n6971), .Y(n4515) );
  AOI22X1 U3788 ( .A(n8924), .B(recentVBools_len_new_reg_317[19]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[19]), .D(n8656), .Y(n2823)
         );
  OAI21X1 U3790 ( .A(ap_CS_fsm[7]), .B(n10127), .C(n7884), .Y(n4516) );
  AOI22X1 U3791 ( .A(n8924), .B(recentVBools_len_new_reg_317[18]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[18]), .D(n8656), .Y(n2825)
         );
  OAI21X1 U3792 ( .A(ap_CS_fsm[7]), .B(n10126), .C(n6369), .Y(n4517) );
  AOI22X1 U3793 ( .A(n8924), .B(recentVBools_len_new_reg_317[17]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[17]), .D(n8656), .Y(n2827)
         );
  OAI21X1 U3794 ( .A(ap_CS_fsm[7]), .B(n10125), .C(n6270), .Y(n4518) );
  AOI22X1 U3795 ( .A(n8924), .B(recentVBools_len_new_reg_317[16]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[16]), .D(n8656), .Y(n2829)
         );
  OAI21X1 U3796 ( .A(ap_CS_fsm[7]), .B(n10124), .C(n6181), .Y(n4519) );
  AOI22X1 U3797 ( .A(n8924), .B(recentVBools_len_new_reg_317[15]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[15]), .D(n8656), .Y(n2831)
         );
  OAI21X1 U3798 ( .A(n9012), .B(n10123), .C(n6108), .Y(n4520) );
  AOI22X1 U3799 ( .A(n8924), .B(recentVBools_len_new_reg_317[14]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[14]), .D(n8656), .Y(n2833)
         );
  OAI21X1 U3800 ( .A(n9012), .B(n10122), .C(n6048), .Y(n4521) );
  AOI22X1 U3801 ( .A(n8924), .B(recentVBools_len_new_reg_317[13]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[13]), .D(n8656), .Y(n2835)
         );
  OAI21X1 U3802 ( .A(ap_CS_fsm[7]), .B(n10121), .C(n7120), .Y(n4522) );
  AOI22X1 U3803 ( .A(n8924), .B(recentVBools_len_new_reg_317[12]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[12]), .D(n8656), .Y(n2837)
         );
  OAI21X1 U3804 ( .A(n9012), .B(n10120), .C(n6969), .Y(n4523) );
  AOI22X1 U3805 ( .A(n8924), .B(recentVBools_len_new_reg_317[11]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[11]), .D(n8656), .Y(n2839)
         );
  OAI21X1 U3806 ( .A(n9012), .B(n10119), .C(n6830), .Y(n4524) );
  AOI22X1 U3807 ( .A(n8924), .B(recentVBools_len_new_reg_317[10]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[10]), .D(n8656), .Y(n2841)
         );
  OAI21X1 U3809 ( .A(ap_CS_fsm[7]), .B(n10118), .C(n6702), .Y(n4525) );
  AOI22X1 U3810 ( .A(n8924), .B(recentVBools_len_new_reg_317[9]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[9]), .D(n8656), .Y(n2843)
         );
  OAI21X1 U3812 ( .A(n9012), .B(n10117), .C(n6586), .Y(n4526) );
  AOI22X1 U3813 ( .A(n8924), .B(recentVBools_len_new_reg_317[8]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[8]), .D(n8656), .Y(n2845)
         );
  OAI21X1 U3815 ( .A(n9012), .B(n10116), .C(n6476), .Y(n4527) );
  AOI22X1 U3816 ( .A(n8924), .B(recentVBools_len_new_reg_317[7]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[7]), .D(n8656), .Y(n2847)
         );
  OAI21X1 U3817 ( .A(ap_CS_fsm[7]), .B(n10115), .C(n8135), .Y(n4528) );
  AOI22X1 U3818 ( .A(n8924), .B(recentVBools_len_new_reg_317[6]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[6]), .D(n8656), .Y(n2849)
         );
  OAI21X1 U3819 ( .A(ap_CS_fsm[7]), .B(n10114), .C(n6368), .Y(n4529) );
  AOI22X1 U3820 ( .A(n8924), .B(recentVBools_len_new_reg_317[5]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[5]), .D(n8656), .Y(n2851)
         );
  OAI21X1 U3821 ( .A(ap_CS_fsm[7]), .B(n10113), .C(n6268), .Y(n4530) );
  AOI22X1 U3822 ( .A(n8924), .B(recentVBools_len_new_reg_317[4]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[4]), .D(n8656), .Y(n2853)
         );
  OAI21X1 U3823 ( .A(ap_CS_fsm[7]), .B(n10112), .C(n6180), .Y(n4531) );
  AOI22X1 U3824 ( .A(n8924), .B(recentVBools_len_new_reg_317[3]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[3]), .D(n8656), .Y(n2855)
         );
  OAI21X1 U3825 ( .A(ap_CS_fsm[7]), .B(n10111), .C(n6107), .Y(n4532) );
  AOI22X1 U3826 ( .A(n8924), .B(recentVBools_len_new_reg_317[2]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[2]), .D(n8656), .Y(n2857)
         );
  OAI21X1 U3828 ( .A(n9012), .B(n10110), .C(n6047), .Y(n4533) );
  AOI22X1 U3829 ( .A(n8924), .B(recentVBools_len_new_reg_317[1]), .C(n10079), 
        .D(n8656), .Y(n2859) );
  OAI21X1 U3831 ( .A(n9012), .B(n10075), .C(n4796), .Y(n4534) );
  AOI22X1 U3832 ( .A(n8924), .B(recentVBools_len_new_reg_317[0]), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[0]), .D(n8656), .Y(n2861)
         );
  OAI21X1 U3835 ( .A(n7094), .B(n2699), .C(n4795), .Y(n4535) );
  AOI22X1 U3836 ( .A(recentVBools_len_new_reg_317[31]), .B(n2701), .C(
        CircularBuffer_len_write_assig_1_fu_924_p2[31]), .D(n2864), .Y(n2863)
         );
  OAI21X1 U3842 ( .A(n8945), .B(n9792), .C(n8126), .Y(n4536) );
  OAI21X1 U3845 ( .A(n8945), .B(n9791), .C(n7876), .Y(n4537) );
  OAI21X1 U3848 ( .A(n8945), .B(n9790), .C(n7661), .Y(n4538) );
  AOI22X1 U3853 ( .A(VCaptureThresh[31]), .B(n8923), .C(v_length[31]), .D(
        n8940), .Y(n2870) );
  AOI22X1 U3856 ( .A(VCaptureThresh[30]), .B(n8923), .C(v_length[30]), .D(
        n8940), .Y(n2873) );
  AOI22X1 U3859 ( .A(VCaptureThresh[29]), .B(n8923), .C(v_length[29]), .D(
        n8940), .Y(n2875) );
  AOI22X1 U3862 ( .A(VCaptureThresh[28]), .B(n8923), .C(v_length[28]), .D(
        n8940), .Y(n2877) );
  AOI22X1 U3865 ( .A(VCaptureThresh[27]), .B(n8923), .C(v_length[27]), .D(
        n8939), .Y(n2879) );
  AOI22X1 U3868 ( .A(VCaptureThresh[26]), .B(n8923), .C(v_length[26]), .D(
        n8939), .Y(n2881) );
  AOI22X1 U3871 ( .A(VCaptureThresh[25]), .B(n8923), .C(v_length[25]), .D(
        n8939), .Y(n2883) );
  AOI22X1 U3874 ( .A(VCaptureThresh[24]), .B(n8923), .C(v_length[24]), .D(
        n8939), .Y(n2885) );
  AOI22X1 U3877 ( .A(VCaptureThresh[23]), .B(n8923), .C(v_length[23]), .D(
        n8939), .Y(n2887) );
  AOI22X1 U3880 ( .A(VCaptureThresh[22]), .B(n8923), .C(v_length[22]), .D(
        n8939), .Y(n2889) );
  AOI22X1 U3883 ( .A(VCaptureThresh[21]), .B(n8923), .C(v_length[21]), .D(
        n8939), .Y(n2891) );
  AOI22X1 U3886 ( .A(VCaptureThresh[20]), .B(n8923), .C(v_length[20]), .D(
        n8939), .Y(n2893) );
  AOI22X1 U3889 ( .A(VCaptureThresh[19]), .B(n8923), .C(v_length[19]), .D(
        n8939), .Y(n2895) );
  AOI22X1 U3892 ( .A(VCaptureThresh[18]), .B(n8923), .C(v_length[18]), .D(
        n8939), .Y(n2897) );
  AOI22X1 U3895 ( .A(VCaptureThresh[17]), .B(n8923), .C(v_length[17]), .D(
        n8939), .Y(n2899) );
  AOI22X1 U3898 ( .A(VCaptureThresh[16]), .B(n8923), .C(v_length[16]), .D(
        n8939), .Y(n2901) );
  AOI22X1 U3901 ( .A(VCaptureThresh[15]), .B(n8923), .C(v_length[15]), .D(
        n8655), .Y(n2903) );
  AOI22X1 U3904 ( .A(VCaptureThresh[14]), .B(n8923), .C(v_length[14]), .D(
        n8655), .Y(n2905) );
  AOI22X1 U3907 ( .A(VCaptureThresh[13]), .B(n8923), .C(v_length[13]), .D(
        n8655), .Y(n2907) );
  AOI22X1 U3910 ( .A(VCaptureThresh[12]), .B(n8923), .C(v_length[12]), .D(
        n8655), .Y(n2909) );
  AOI22X1 U3913 ( .A(VCaptureThresh[11]), .B(n8923), .C(v_length[11]), .D(
        n8655), .Y(n2911) );
  AOI22X1 U3916 ( .A(VCaptureThresh[10]), .B(n8923), .C(v_length[10]), .D(
        n8655), .Y(n2913) );
  AOI22X1 U3919 ( .A(VCaptureThresh[9]), .B(n8923), .C(v_length[9]), .D(n8655), 
        .Y(n2915) );
  AOI22X1 U3922 ( .A(VCaptureThresh[8]), .B(n8923), .C(v_length[8]), .D(n8655), 
        .Y(n2917) );
  AOI22X1 U3925 ( .A(VCaptureThresh[7]), .B(n8923), .C(v_length[7]), .D(n8936), 
        .Y(n2919) );
  AOI22X1 U3928 ( .A(VCaptureThresh[6]), .B(n8923), .C(v_length[6]), .D(n8936), 
        .Y(n2921) );
  AOI22X1 U3931 ( .A(VCaptureThresh[5]), .B(n8923), .C(v_length[5]), .D(n8936), 
        .Y(n2923) );
  AOI22X1 U3934 ( .A(VCaptureThresh[4]), .B(n8923), .C(v_length[4]), .D(n8936), 
        .Y(n2925) );
  AOI22X1 U3937 ( .A(VCaptureThresh[3]), .B(n8923), .C(v_length[3]), .D(n8936), 
        .Y(n2927) );
  AOI22X1 U3940 ( .A(VCaptureThresh[2]), .B(n8923), .C(v_length[2]), .D(n8936), 
        .Y(n2929) );
  AOI22X1 U3943 ( .A(VCaptureThresh[1]), .B(n8923), .C(v_length[1]), .D(n8936), 
        .Y(n2931) );
  AOI22X1 U3946 ( .A(VCaptureThresh[0]), .B(n8923), .C(v_length[0]), .D(n8936), 
        .Y(n2933) );
  OAI21X1 U3947 ( .A(n8945), .B(n9762), .C(n7454), .Y(n4571) );
  OAI21X1 U3950 ( .A(n8945), .B(n9756), .C(n7274), .Y(n4572) );
  OAI21X1 U3953 ( .A(n8945), .B(n9754), .C(n7108), .Y(n4573) );
  OAI21X1 U3956 ( .A(n8945), .B(n9752), .C(n6957), .Y(n4574) );
  OAI21X1 U3959 ( .A(n8945), .B(n9748), .C(n6818), .Y(n4575) );
  OAI21X1 U3962 ( .A(n8945), .B(n9742), .C(n6693), .Y(n4576) );
  OAI21X1 U3965 ( .A(n8945), .B(n9739), .C(n6578), .Y(n4577) );
  OAI21X1 U3968 ( .A(n8946), .B(n9735), .C(n8125), .Y(n4578) );
  OAI21X1 U3971 ( .A(n8946), .B(n9731), .C(n7875), .Y(n4579) );
  OAI21X1 U3974 ( .A(n8946), .B(n9725), .C(n7660), .Y(n4580) );
  OAI21X1 U3977 ( .A(n8946), .B(n9722), .C(n7453), .Y(n4581) );
  OAI21X1 U3980 ( .A(n8946), .B(n9718), .C(n7273), .Y(n4582) );
  OAI21X1 U3983 ( .A(n8946), .B(n9714), .C(n7107), .Y(n4583) );
  OAI21X1 U3986 ( .A(n8946), .B(n9708), .C(n6956), .Y(n4584) );
  OAI21X1 U3989 ( .A(n8946), .B(n9706), .C(n6817), .Y(n4585) );
  OAI21X1 U3992 ( .A(n8946), .B(n9704), .C(n6692), .Y(n4586) );
  OAI21X1 U3995 ( .A(n8946), .B(n9700), .C(n6577), .Y(n4587) );
  OAI21X1 U3998 ( .A(n8946), .B(n9694), .C(n6464), .Y(n4588) );
  OAI21X1 U4001 ( .A(n8947), .B(n9691), .C(n6463), .Y(n4589) );
  OAI21X1 U4004 ( .A(n8947), .B(n9688), .C(n6355), .Y(n4590) );
  OAI21X1 U4007 ( .A(n8947), .B(n9684), .C(n6259), .Y(n4591) );
  OAI21X1 U4010 ( .A(n8946), .B(n9678), .C(n6170), .Y(n4592) );
  OAI21X1 U4013 ( .A(n8947), .B(n9674), .C(n6098), .Y(n4593) );
  OAI21X1 U4016 ( .A(n8948), .B(n9669), .C(n8124), .Y(n4594) );
  OAI21X1 U4019 ( .A(n8948), .B(n9666), .C(n7874), .Y(n4595) );
  OAI21X1 U4022 ( .A(n8947), .B(n9662), .C(n7659), .Y(n4596) );
  OAI21X1 U4025 ( .A(n8949), .B(n9660), .C(n6258), .Y(n4597) );
  OAI21X1 U4028 ( .A(n8947), .B(n9658), .C(n6169), .Y(n4598) );
  OAI21X1 U4031 ( .A(n8949), .B(n9655), .C(n6462), .Y(n4599) );
  OAI21X1 U4034 ( .A(n8948), .B(n9651), .C(n6354), .Y(n4600) );
  OAI21X1 U4037 ( .A(n8949), .B(n9648), .C(n6038), .Y(n4601) );
  OAI21X1 U4040 ( .A(n8949), .B(n9647), .C(n6097), .Y(n4602) );
  AOI22X1 U4045 ( .A(ACaptureThresh[31]), .B(n8923), .C(a_length[31]), .D(
        n8936), .Y(n2999) );
  AOI22X1 U4048 ( .A(ACaptureThresh[30]), .B(n8923), .C(a_length[30]), .D(
        n8936), .Y(n3001) );
  AOI22X1 U4051 ( .A(ACaptureThresh[29]), .B(n8923), .C(a_length[29]), .D(
        n8936), .Y(n3003) );
  AOI22X1 U4054 ( .A(ACaptureThresh[28]), .B(n8923), .C(a_length[28]), .D(
        n8936), .Y(n3005) );
  AOI22X1 U4057 ( .A(ACaptureThresh[27]), .B(n8923), .C(a_length[27]), .D(
        n8937), .Y(n3007) );
  AOI22X1 U4060 ( .A(ACaptureThresh[26]), .B(n8923), .C(a_length[26]), .D(
        n8937), .Y(n3009) );
  AOI22X1 U4063 ( .A(ACaptureThresh[25]), .B(n8923), .C(a_length[25]), .D(
        n8937), .Y(n3011) );
  AOI22X1 U4066 ( .A(ACaptureThresh[24]), .B(n8923), .C(a_length[24]), .D(
        n8937), .Y(n3013) );
  AOI22X1 U4069 ( .A(ACaptureThresh[23]), .B(n8923), .C(a_length[23]), .D(
        n8937), .Y(n3015) );
  AOI22X1 U4072 ( .A(ACaptureThresh[22]), .B(n8923), .C(a_length[22]), .D(
        n8937), .Y(n3017) );
  AOI22X1 U4075 ( .A(ACaptureThresh[21]), .B(n8923), .C(a_length[21]), .D(
        n8937), .Y(n3019) );
  AOI22X1 U4078 ( .A(ACaptureThresh[20]), .B(n8923), .C(a_length[20]), .D(
        n8937), .Y(n3021) );
  AOI22X1 U4081 ( .A(ACaptureThresh[19]), .B(n8923), .C(a_length[19]), .D(
        n8937), .Y(n3023) );
  AOI22X1 U4084 ( .A(ACaptureThresh[18]), .B(n8923), .C(a_length[18]), .D(
        n8937), .Y(n3025) );
  AOI22X1 U4087 ( .A(ACaptureThresh[17]), .B(n8923), .C(a_length[17]), .D(
        n8937), .Y(n3027) );
  AOI22X1 U4090 ( .A(ACaptureThresh[16]), .B(n8923), .C(a_length[16]), .D(
        n8937), .Y(n3029) );
  AOI22X1 U4093 ( .A(ACaptureThresh[15]), .B(n8923), .C(a_length[15]), .D(
        n8938), .Y(n3031) );
  AOI22X1 U4096 ( .A(ACaptureThresh[14]), .B(n8923), .C(a_length[14]), .D(
        n8938), .Y(n3033) );
  AOI22X1 U4099 ( .A(ACaptureThresh[13]), .B(n8923), .C(a_length[13]), .D(
        n8938), .Y(n3035) );
  AOI22X1 U4102 ( .A(ACaptureThresh[12]), .B(n8923), .C(a_length[12]), .D(
        n8938), .Y(n3037) );
  AOI22X1 U4105 ( .A(ACaptureThresh[11]), .B(n8923), .C(a_length[11]), .D(
        n8938), .Y(n3039) );
  AOI22X1 U4108 ( .A(ACaptureThresh[10]), .B(n8923), .C(a_length[10]), .D(
        n8938), .Y(n3041) );
  AOI22X1 U4111 ( .A(ACaptureThresh[9]), .B(n8923), .C(a_length[9]), .D(n8938), 
        .Y(n3043) );
  AOI22X1 U4114 ( .A(ACaptureThresh[8]), .B(n8923), .C(a_length[8]), .D(n8938), 
        .Y(n3045) );
  AOI22X1 U4117 ( .A(ACaptureThresh[7]), .B(n8923), .C(a_length[7]), .D(n8938), 
        .Y(n3047) );
  AOI22X1 U4120 ( .A(ACaptureThresh[6]), .B(n8923), .C(a_length[6]), .D(n8938), 
        .Y(n3049) );
  AOI22X1 U4123 ( .A(ACaptureThresh[5]), .B(n8923), .C(a_length[5]), .D(n8938), 
        .Y(n3051) );
  AOI22X1 U4126 ( .A(ACaptureThresh[4]), .B(n8923), .C(a_length[4]), .D(n8938), 
        .Y(n3053) );
  AOI22X1 U4129 ( .A(ACaptureThresh[3]), .B(n8923), .C(a_length[3]), .D(n8939), 
        .Y(n3055) );
  AOI22X1 U4132 ( .A(ACaptureThresh[2]), .B(n8923), .C(a_length[2]), .D(n8936), 
        .Y(n3057) );
  AOI22X1 U4135 ( .A(ACaptureThresh[1]), .B(n8923), .C(a_length[1]), .D(n8655), 
        .Y(n3059) );
  AOI22X1 U4138 ( .A(ACaptureThresh[0]), .B(n8923), .C(a_length[0]), .D(n8655), 
        .Y(n3061) );
  OAI21X1 U4140 ( .A(n8949), .B(n9645), .C(n5050), .Y(n4635) );
  OAI21X1 U4143 ( .A(n8949), .B(n9639), .C(n5049), .Y(n4636) );
  OAI21X1 U4146 ( .A(n8948), .B(n9637), .C(n7452), .Y(n4637) );
  OAI21X1 U4149 ( .A(n8949), .B(n9635), .C(n7272), .Y(n4638) );
  OAI21X1 U4152 ( .A(n8950), .B(n9633), .C(n7106), .Y(n4639) );
  OAI21X1 U4155 ( .A(n8950), .B(n9627), .C(n6955), .Y(n4640) );
  OAI21X1 U4158 ( .A(n8949), .B(n9625), .C(n6816), .Y(n4641) );
  OAI21X1 U4161 ( .A(n8950), .B(n9621), .C(n6691), .Y(n4642) );
  OAI21X1 U4164 ( .A(n8950), .B(n9619), .C(n6576), .Y(n4643) );
  OAI21X1 U4167 ( .A(n8948), .B(n9613), .C(n6461), .Y(n4644) );
  OAI21X1 U4170 ( .A(n8950), .B(n9611), .C(n6353), .Y(n4645) );
  OAI21X1 U4173 ( .A(n8948), .B(n9607), .C(n6257), .Y(n4646) );
  OAI21X1 U4176 ( .A(n8950), .B(n9605), .C(n6168), .Y(n4647) );
  OAI21X1 U4179 ( .A(n8951), .B(n9599), .C(n6096), .Y(n4648) );
  OAI21X1 U4182 ( .A(n8951), .B(n9597), .C(n6037), .Y(n4649) );
  OAI21X1 U4185 ( .A(n8950), .B(n9595), .C(n5048), .Y(n4650) );
  OAI21X1 U4188 ( .A(n8951), .B(n9593), .C(n5047), .Y(n4651) );
  OAI21X1 U4191 ( .A(n8951), .B(n9587), .C(n8123), .Y(n4652) );
  OAI21X1 U4194 ( .A(n8947), .B(n9585), .C(n7873), .Y(n4653) );
  OAI21X1 U4197 ( .A(n8950), .B(n9582), .C(n7658), .Y(n4654) );
  OAI21X1 U4200 ( .A(n8950), .B(n9580), .C(n7451), .Y(n4655) );
  OAI21X1 U4203 ( .A(n8951), .B(n9574), .C(n7271), .Y(n4656) );
  OAI21X1 U4206 ( .A(n8950), .B(n9572), .C(n6815), .Y(n4657) );
  OAI21X1 U4209 ( .A(n8950), .B(n9567), .C(n6256), .Y(n4658) );
  OAI21X1 U4212 ( .A(n8950), .B(n9565), .C(n6095), .Y(n4659) );
  OAI21X1 U4215 ( .A(n8949), .B(n9561), .C(n6954), .Y(n4660) );
  OAI21X1 U4218 ( .A(n8949), .B(n9559), .C(n7105), .Y(n4661) );
  OAI21X1 U4221 ( .A(n8950), .B(n9557), .C(n6036), .Y(n4662) );
  OAI21X1 U4224 ( .A(n8949), .B(n9555), .C(n6690), .Y(n4663) );
  OAI21X1 U4227 ( .A(n8949), .B(n9551), .C(n6575), .Y(n4664) );
  OAI21X1 U4230 ( .A(n8949), .B(n9549), .C(n7872), .Y(n4665) );
  OAI21X1 U4233 ( .A(n8948), .B(n9548), .C(n7657), .Y(n4666) );
  OAI21X1 U4236 ( .A(n8948), .B(n9547), .C(n7104), .Y(n4667) );
  OAI21X1 U4239 ( .A(n8948), .B(n9546), .C(n6953), .Y(n4668) );
  OAI21X1 U4242 ( .A(n8947), .B(n9545), .C(n6814), .Y(n4669) );
  OAI21X1 U4245 ( .A(n8948), .B(n9544), .C(n6167), .Y(n4670) );
  OAI21X1 U4248 ( .A(n8948), .B(n9543), .C(n5046), .Y(n4671) );
  OAI21X1 U4251 ( .A(n8948), .B(n9542), .C(n5045), .Y(n4672) );
  OAI21X1 U4254 ( .A(n8948), .B(n9541), .C(n6689), .Y(n4673) );
  OAI21X1 U4257 ( .A(n8947), .B(n9533), .C(n7450), .Y(n4674) );
  OAI21X1 U4260 ( .A(n8947), .B(n9495), .C(n6574), .Y(n4675) );
  OAI21X1 U4263 ( .A(n8947), .B(n9494), .C(n5044), .Y(n4676) );
  OAI21X1 U4266 ( .A(n8946), .B(n9493), .C(n6352), .Y(n4677) );
  OAI21X1 U4269 ( .A(n8947), .B(n9492), .C(n5043), .Y(n4678) );
  OAI21X1 U4272 ( .A(n8947), .B(n9491), .C(n5042), .Y(n4679) );
  OAI21X1 U4277 ( .A(n10740), .B(n2202), .C(n8173), .Y(n4680) );
  OAI21X1 U4280 ( .A(\last_sample_is_A_V[0] ), .B(n5966), .C(ap_CS_fsm[12]), 
        .Y(n2202) );
  NAND3X1 U4281 ( .A(N499), .B(N498), .C(n5876), .Y(n2237) );
  NAND3X1 U4285 ( .A(n8304), .B(n10670), .C(ap_rst_n), .Y(N98) );
  AOI21X1 U4307 ( .A(n10535), .B(n8934), .C(n9042), .Y(N110) );
  AOI21X1 U4317 ( .A(n10057), .B(n8927), .C(n9042), .Y(N105) );
  OAI21X1 U4449 ( .A(n8920), .B(n10217), .C(n6784), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[9]) );
  OAI21X1 U4452 ( .A(n8920), .B(n10216), .C(n6919), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[8]) );
  OAI21X1 U4455 ( .A(n8920), .B(n10215), .C(n7061), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[7]) );
  OAI21X1 U4458 ( .A(n8920), .B(n10214), .C(n7215), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[6]) );
  OAI21X1 U4461 ( .A(n8920), .B(n10213), .C(n7373), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[5]) );
  OAI21X1 U4464 ( .A(n8920), .B(n10212), .C(n7556), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[4]) );
  OAI21X1 U4467 ( .A(n8920), .B(n10211), .C(n7755), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[3]) );
  OAI21X1 U4470 ( .A(n8920), .B(n10241), .C(n8216), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[31]) );
  OAI21X1 U4473 ( .A(n8920), .B(n10238), .C(n6233), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[30]) );
  OAI21X1 U4476 ( .A(n8920), .B(n10210), .C(n7970), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[2]) );
  OAI21X1 U4479 ( .A(n8920), .B(n10237), .C(n5041), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[29]) );
  OAI21X1 U4482 ( .A(n8920), .B(n10236), .C(n6551), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[28]) );
  OAI21X1 U4485 ( .A(n8920), .B(n10235), .C(n6780), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[27]) );
  OAI21X1 U4488 ( .A(n8920), .B(n10234), .C(n5040), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[26]) );
  OAI21X1 U4491 ( .A(n8920), .B(n10233), .C(n5039), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[25]) );
  OAI21X1 U4494 ( .A(n8920), .B(n10232), .C(n6153), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[24]) );
  OAI21X1 U4497 ( .A(n8920), .B(n10231), .C(n6238), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[23]) );
  OAI21X1 U4500 ( .A(n8920), .B(n10230), .C(n6331), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[22]) );
  OAI21X1 U4503 ( .A(n8920), .B(n10229), .C(n6440), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[21]) );
  OAI21X1 U4506 ( .A(n8920), .B(n10228), .C(n6662), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[20]) );
  OAI21X1 U4509 ( .A(n8920), .B(n10209), .C(n8211), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[1]) );
  OAI21X1 U4512 ( .A(n8920), .B(n10227), .C(n6917), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[19]) );
  OAI21X1 U4515 ( .A(n8920), .B(n10226), .C(n7059), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[18]) );
  OAI21X1 U4518 ( .A(n8920), .B(n10225), .C(n6333), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[17]) );
  OAI21X1 U4521 ( .A(n8920), .B(n10224), .C(n7213), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[16]) );
  OAI21X1 U4524 ( .A(n8920), .B(n10223), .C(n7371), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[15]) );
  OAI21X1 U4527 ( .A(n8920), .B(n10222), .C(n7554), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[14]) );
  OAI21X1 U4530 ( .A(n8920), .B(n10221), .C(n7753), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[13]) );
  OAI21X1 U4533 ( .A(n8920), .B(n10220), .C(n6442), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[12]) );
  OAI21X1 U4536 ( .A(n8920), .B(n10219), .C(n6553), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[11]) );
  OAI21X1 U4539 ( .A(n8920), .B(n10218), .C(n6664), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[10]) );
  OAI21X1 U4542 ( .A(n8920), .B(n10208), .C(n7972), .Y(
        CircularBuffer_int_30_sum_i_fu_758_p3[0]) );
  NAND3X1 U4547 ( .A(n3187), .B(n3188), .C(n3189), .Y(n3186) );
  NOR3X1 U4548 ( .A(n7821), .B(n7819), .C(n7820), .Y(n3189) );
  NAND3X1 U4555 ( .A(n10126), .B(n10127), .C(n8260), .Y(n3190) );
  NOR3X1 U4559 ( .A(n7416), .B(recentVBools_len[10]), .C(recentVBools_len[0]), 
        .Y(n3188) );
  NOR3X1 U4563 ( .A(n7240), .B(n10112), .C(n10113), .Y(n3187) );
  NAND3X1 U4567 ( .A(n3196), .B(n3197), .C(n3198), .Y(n3185) );
  NOR3X1 U4568 ( .A(n8034), .B(n8032), .C(n8033), .Y(n3198) );
  NAND3X1 U4575 ( .A(n10115), .B(n10116), .C(n8261), .Y(n3199) );
  NOR3X1 U4579 ( .A(n8283), .B(recentVBools_len[26]), .C(recentVBools_len[25]), 
        .Y(n3197) );
  NOR3X1 U4583 ( .A(n7603), .B(recentVBools_len[22]), .C(recentVBools_len[21]), 
        .Y(n3196) );
  OAI21X1 U4587 ( .A(n8922), .B(n10552), .C(n6785), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[9]) );
  OAI21X1 U4590 ( .A(n8922), .B(n10551), .C(n6920), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[8]) );
  OAI21X1 U4593 ( .A(n8922), .B(n10550), .C(n7062), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[7]) );
  OAI21X1 U4596 ( .A(n8922), .B(n10549), .C(n7216), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[6]) );
  OAI21X1 U4599 ( .A(n8922), .B(n10548), .C(n7374), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[5]) );
  OAI21X1 U4602 ( .A(n8922), .B(n10547), .C(n7557), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[4]) );
  OAI21X1 U4605 ( .A(n8922), .B(n10546), .C(n7756), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[3]) );
  OAI21X1 U4608 ( .A(n8922), .B(n9384), .C(n8217), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[31]) );
  OAI21X1 U4611 ( .A(n8922), .B(n10811), .C(n6234), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[30]) );
  OAI21X1 U4614 ( .A(n8922), .B(n10545), .C(n7971), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[2]) );
  OAI21X1 U4617 ( .A(n8922), .B(n10572), .C(n5038), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[29]) );
  OAI21X1 U4620 ( .A(n8922), .B(n10571), .C(n6552), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[28]) );
  OAI21X1 U4623 ( .A(n8922), .B(n10570), .C(n6782), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[27]) );
  OAI21X1 U4626 ( .A(n8922), .B(n10569), .C(n5037), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[26]) );
  OAI21X1 U4629 ( .A(n8922), .B(n10568), .C(n5036), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[25]) );
  OAI21X1 U4632 ( .A(n8922), .B(n10567), .C(n6154), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[24]) );
  OAI21X1 U4635 ( .A(n8922), .B(n10566), .C(n6239), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[23]) );
  OAI21X1 U4638 ( .A(n8922), .B(n10565), .C(n6332), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[22]) );
  OAI21X1 U4641 ( .A(n8922), .B(n10564), .C(n6441), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[21]) );
  OAI21X1 U4644 ( .A(n8922), .B(n10563), .C(n6663), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[20]) );
  OAI21X1 U4647 ( .A(n8922), .B(n10544), .C(n8212), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[1]) );
  OAI21X1 U4650 ( .A(n8922), .B(n10562), .C(n6918), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[19]) );
  OAI21X1 U4653 ( .A(n8922), .B(n10561), .C(n7060), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[18]) );
  OAI21X1 U4656 ( .A(n8922), .B(n10560), .C(n6334), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[17]) );
  OAI21X1 U4659 ( .A(n8922), .B(n10559), .C(n7214), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[16]) );
  OAI21X1 U4662 ( .A(n8922), .B(n10558), .C(n7372), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[15]) );
  OAI21X1 U4665 ( .A(n8922), .B(n10557), .C(n7555), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[14]) );
  OAI21X1 U4668 ( .A(n8922), .B(n10556), .C(n7754), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[13]) );
  OAI21X1 U4671 ( .A(n8922), .B(n10555), .C(n6443), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[12]) );
  OAI21X1 U4674 ( .A(n8922), .B(n10554), .C(n6554), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[11]) );
  OAI21X1 U4677 ( .A(n8922), .B(n10553), .C(n6665), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[10]) );
  OAI21X1 U4680 ( .A(n8922), .B(n10543), .C(n7973), .Y(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[0]) );
  NAND3X1 U4685 ( .A(n3239), .B(n3240), .C(n3241), .Y(n3238) );
  NOR3X1 U4686 ( .A(n7824), .B(n7822), .C(n7823), .Y(n3241) );
  NAND3X1 U4693 ( .A(n10621), .B(n10622), .C(n8262), .Y(n3242) );
  NOR3X1 U4697 ( .A(n7417), .B(recentABools_len[10]), .C(recentABools_len[0]), 
        .Y(n3240) );
  NOR3X1 U4701 ( .A(n7241), .B(n10607), .C(n10608), .Y(n3239) );
  NAND3X1 U4705 ( .A(n3248), .B(n3249), .C(n3250), .Y(n3237) );
  NOR3X1 U4706 ( .A(n8037), .B(n8035), .C(n8036), .Y(n3250) );
  NAND3X1 U4713 ( .A(n10610), .B(n10611), .C(n8263), .Y(n3251) );
  NOR3X1 U4717 ( .A(n8284), .B(recentABools_len[26]), .C(recentABools_len[25]), 
        .Y(n3249) );
  NOR3X1 U4721 ( .A(n7604), .B(recentABools_len[22]), .C(recentABools_len[21]), 
        .Y(n3248) );
  AOI21X1 \Decision_AXILiteS_s_axi_U/U879  ( .A(n10884), .B(n10885), .C(n10888), .Y(interrupt) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U878  ( .A(ap_rst_n), .B(n9280), .C(
        s_axi_AXILiteS_WREADY), .Y(\Decision_AXILiteS_s_axi_U/n645 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U877  ( .A(s_axi_AXILiteS_AWREADY), .B(
        ap_rst_n), .C(s_axi_AXILiteS_AWVALID), .Y(
        \Decision_AXILiteS_s_axi_U/n646 ) );
  NOR3X1 \Decision_AXILiteS_s_axi_U/U874  ( .A(n8354), .B(
        s_axi_AXILiteS_BREADY), .C(n9042), .Y(\Decision_AXILiteS_s_axi_U/n644 ) );
  AOI21X1 \Decision_AXILiteS_s_axi_U/U873  ( .A(
        \Decision_AXILiteS_s_axi_U/n625 ), .B(ap_rst_n), .C(
        \Decision_AXILiteS_s_axi_U/n644 ), .Y(\Decision_AXILiteS_s_axi_U/n643 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U869  ( .A(n8652), .B(n10899), .C(n8182), 
        .Y(\Decision_AXILiteS_s_axi_U/n871 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U867  ( .A(n8652), .B(n10898), .C(n7940), 
        .Y(\Decision_AXILiteS_s_axi_U/n870 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U865  ( .A(n8652), .B(n10897), .C(n7723), 
        .Y(\Decision_AXILiteS_s_axi_U/n869 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U863  ( .A(n8652), .B(n10895), .C(n7525), 
        .Y(\Decision_AXILiteS_s_axi_U/n868 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U861  ( .A(n8652), .B(n10894), .C(n7346), 
        .Y(\Decision_AXILiteS_s_axi_U/n867 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U859  ( .A(n8652), .B(n10893), .C(n7183), 
        .Y(\Decision_AXILiteS_s_axi_U/n866 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U857  ( .A(n8652), .B(n10892), .C(n7030), 
        .Y(\Decision_AXILiteS_s_axi_U/n865 ) );
  NOR3X1 \Decision_AXILiteS_s_axi_U/U854  ( .A(s_axi_AXILiteS_ARREADY), .B(
        s_axi_AXILiteS_RREADY), .C(n9042), .Y(\Decision_AXILiteS_s_axi_U/n634 ) );
  AOI21X1 \Decision_AXILiteS_s_axi_U/U853  ( .A(ap_rst_n), .B(
        \Decision_AXILiteS_s_axi_U/n630 ), .C(\Decision_AXILiteS_s_axi_U/n634 ), .Y(\Decision_AXILiteS_s_axi_U/n633 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U850  ( .A(
        \Decision_AXILiteS_s_axi_U/n310 ), .B(n9321), .C(n5894), .Y(
        \Decision_AXILiteS_s_axi_U/n631 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U848  ( .A(ap_rst_n), .B(n9316), .C(n8266), .Y(\Decision_AXILiteS_s_axi_U/n628 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U845  ( .A(
        \Decision_AXILiteS_s_axi_U/int_ap_done ), .B(n5570), .C(n8429), .Y(
        \Decision_AXILiteS_s_axi_U/n626 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U842  ( .A(n10892), .B(n10893), .C(
        \Decision_AXILiteS_s_axi_U/n625 ), .Y(\Decision_AXILiteS_s_axi_U/n616 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U840  ( .A(n10898), .B(n10899), .C(n10897), .Y(\Decision_AXILiteS_s_axi_U/n615 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U839  ( .A(n8382), .B(n10895), .C(n10896), 
        .Y(\Decision_AXILiteS_s_axi_U/n622 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U838  ( .A(n5955), .B(n5964), .C(ap_rst_n), .Y(\Decision_AXILiteS_s_axi_U/n623 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U837  ( .A(ap_rst_n), .B(
        \Decision_AXILiteS_s_axi_U/n623 ), .C(s_axi_AXILiteS_WDATA[7]), .Y(
        \Decision_AXILiteS_s_axi_U/n624 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U836  ( .A(n10890), .B(
        \Decision_AXILiteS_s_axi_U/n623 ), .C(n4926), .Y(
        \Decision_AXILiteS_s_axi_U/n862 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U835  ( .A(
        \Decision_AXILiteS_s_axi_U/int_auto_restart ), .B(ap_CS_fsm[13]), .C(
        \Decision_AXILiteS_s_axi_U/n621 ), .D(n5963), .Y(
        \Decision_AXILiteS_s_axi_U/n618 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U833  ( .A(n5500), .B(ap_rst_n), .C(
        ap_start), .Y(\Decision_AXILiteS_s_axi_U/n619 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U832  ( .A(n5532), .B(n9042), .C(n4925), 
        .Y(\Decision_AXILiteS_s_axi_U/n861 ) );
  NOR3X1 \Decision_AXILiteS_s_axi_U/U831  ( .A(n7631), .B(n7847), .C(n10894), 
        .Y(\Decision_AXILiteS_s_axi_U/n606 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U830  ( .A(
        \Decision_AXILiteS_s_axi_U/n617 ), .B(n10895), .C(
        \Decision_AXILiteS_s_axi_U/n606 ), .Y(\Decision_AXILiteS_s_axi_U/n614 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U828  ( .A(ap_rst_n), .B(n6009), .C(
        s_axi_AXILiteS_WDATA[0]), .Y(\Decision_AXILiteS_s_axi_U/n613 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U827  ( .A(n10888), .B(n6009), .C(n4924), 
        .Y(\Decision_AXILiteS_s_axi_U/n860 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U826  ( .A(
        \Decision_AXILiteS_s_axi_U/n617 ), .B(n8382), .C(
        \Decision_AXILiteS_s_axi_U/n611 ), .Y(\Decision_AXILiteS_s_axi_U/n610 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U824  ( .A(ap_rst_n), .B(n8105), .C(
        s_axi_AXILiteS_WDATA[1]), .Y(\Decision_AXILiteS_s_axi_U/n609 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U823  ( .A(n10887), .B(n8105), .C(n4923), 
        .Y(\Decision_AXILiteS_s_axi_U/n859 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U822  ( .A(ap_rst_n), .B(n8105), .C(
        s_axi_AXILiteS_WDATA[0]), .Y(\Decision_AXILiteS_s_axi_U/n608 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U821  ( .A(n10886), .B(n8105), .C(n4922), 
        .Y(\Decision_AXILiteS_s_axi_U/n858 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U820  ( .A(
        \Decision_AXILiteS_s_axi_U/waddr[3] ), .B(s_axi_AXILiteS_WSTRB[0]), 
        .C(\Decision_AXILiteS_s_axi_U/n606 ), .Y(
        \Decision_AXILiteS_s_axi_U/n605 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U817  ( .A(n8388), .B(
        s_axi_AXILiteS_WDATA[0]), .C(n7625), .Y(
        \Decision_AXILiteS_s_axi_U/n604 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U816  ( .A(s_axi_AXILiteS_WDATA[0]), .B(
        n10885), .C(n9281), .Y(\Decision_AXILiteS_s_axi_U/n603 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U815  ( .A(n10886), .B(n10670), .C(n4921), 
        .Y(\Decision_AXILiteS_s_axi_U/n602 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U813  ( .A(n9277), .B(n10885), .C(n7375), 
        .Y(\Decision_AXILiteS_s_axi_U/n857 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U812  ( .A(s_axi_AXILiteS_WDATA[1]), .B(
        n10884), .C(\Decision_AXILiteS_s_axi_U/n599 ), .Y(
        \Decision_AXILiteS_s_axi_U/n595 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U811  ( .A(
        \Decision_AXILiteS_s_axi_U/int_ier[1] ), .B(ap_CS_fsm[13]), .C(
        ap_rst_n), .Y(\Decision_AXILiteS_s_axi_U/n596 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U810  ( .A(s_axi_AXILiteS_WDATA[1]), .B(
        n8388), .C(n7625), .Y(\Decision_AXILiteS_s_axi_U/n598 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U808  ( .A(n5483), .B(n5569), .C(n5893), 
        .Y(\Decision_AXILiteS_s_axi_U/n856 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U806  ( .A(n10883), .B(n8883), .C(n5035), 
        .Y(\Decision_AXILiteS_s_axi_U/n855 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U804  ( .A(n10882), .B(n8883), .C(n5035), 
        .Y(\Decision_AXILiteS_s_axi_U/n854 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U802  ( .A(n10881), .B(n8883), .C(n5035), 
        .Y(\Decision_AXILiteS_s_axi_U/n853 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U800  ( .A(n10880), .B(n8883), .C(n5035), 
        .Y(\Decision_AXILiteS_s_axi_U/n852 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U798  ( .A(n10879), .B(n8883), .C(n5034), 
        .Y(\Decision_AXILiteS_s_axi_U/n851 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U796  ( .A(n10878), .B(n8883), .C(n5034), 
        .Y(\Decision_AXILiteS_s_axi_U/n850 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U794  ( .A(n10877), .B(n8883), .C(n5034), 
        .Y(\Decision_AXILiteS_s_axi_U/n849 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U792  ( .A(n10876), .B(n8883), .C(n5034), 
        .Y(\Decision_AXILiteS_s_axi_U/n848 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U790  ( .A(n10875), .B(n8883), .C(n6763), 
        .Y(\Decision_AXILiteS_s_axi_U/n847 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U788  ( .A(n10874), .B(n8883), .C(n6763), 
        .Y(\Decision_AXILiteS_s_axi_U/n846 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U786  ( .A(n10873), .B(n8883), .C(n6763), 
        .Y(\Decision_AXILiteS_s_axi_U/n845 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U784  ( .A(n10872), .B(n8883), .C(n6763), 
        .Y(\Decision_AXILiteS_s_axi_U/n844 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U782  ( .A(n10871), .B(n8883), .C(n5033), 
        .Y(\Decision_AXILiteS_s_axi_U/n843 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U780  ( .A(n10870), .B(n8883), .C(n5033), 
        .Y(\Decision_AXILiteS_s_axi_U/n842 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U778  ( .A(n10869), .B(n8883), .C(n5033), 
        .Y(\Decision_AXILiteS_s_axi_U/n841 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U776  ( .A(n10868), .B(n8883), .C(n5033), 
        .Y(\Decision_AXILiteS_s_axi_U/n840 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U774  ( .A(
        \Decision_AXILiteS_s_axi_U/n417 ), .B(\Decision_AXILiteS_s_axi_U/n371 ), .C(\Decision_AXILiteS_s_axi_U/n575 ), .Y(\Decision_AXILiteS_s_axi_U/n574 )
         );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U771  ( .A(n8104), .B(
        \Decision_AXILiteS_s_axi_U/n572 ), .C(\reset_A_V[0] ), .Y(
        \Decision_AXILiteS_s_axi_U/n573 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U770  ( .A(
        \Decision_AXILiteS_s_axi_U/n572 ), .B(n8389), .C(
        \Decision_AXILiteS_s_axi_U/n573 ), .Y(\Decision_AXILiteS_s_axi_U/n839 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U768  ( .A(
        \Decision_AXILiteS_s_axi_U/n371 ), .B(n10899), .C(
        \Decision_AXILiteS_s_axi_U/waddr[5] ), .Y(
        \Decision_AXILiteS_s_axi_U/n522 ) );
  AOI21X1 \Decision_AXILiteS_s_axi_U/U767  ( .A(
        \Decision_AXILiteS_s_axi_U/n481 ), .B(n9278), .C(n9042), .Y(
        \Decision_AXILiteS_s_axi_U/n570 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U766  ( .A(n8104), .B(n7855), .C(
        \reset_V_V[0] ), .Y(\Decision_AXILiteS_s_axi_U/n571 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U765  ( .A(n7855), .B(n8389), .C(
        \Decision_AXILiteS_s_axi_U/n571 ), .Y(\Decision_AXILiteS_s_axi_U/n838 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U764  ( .A(
        \Decision_AXILiteS_s_axi_U/waddr[3] ), .B(n10897), .C(n9278), .Y(
        \Decision_AXILiteS_s_axi_U/n569 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U763  ( .A(n8104), .B(
        \Decision_AXILiteS_s_axi_U/n567 ), .C(\reset_params_V[0] ), .Y(
        \Decision_AXILiteS_s_axi_U/n568 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U762  ( .A(
        \Decision_AXILiteS_s_axi_U/n567 ), .B(n8389), .C(
        \Decision_AXILiteS_s_axi_U/n568 ), .Y(\Decision_AXILiteS_s_axi_U/n837 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U761  ( .A(
        \Decision_AXILiteS_s_axi_U/waddr[4] ), .B(n10895), .C(n9278), .Y(
        \Decision_AXILiteS_s_axi_U/n566 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U758  ( .A(
        \Decision_AXILiteS_s_axi_U/n555 ), .B(n10860), .C(n6217), .Y(
        \Decision_AXILiteS_s_axi_U/n836 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U756  ( .A(
        \Decision_AXILiteS_s_axi_U/n555 ), .B(n10861), .C(n6311), .Y(
        \Decision_AXILiteS_s_axi_U/n835 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U754  ( .A(
        \Decision_AXILiteS_s_axi_U/n555 ), .B(n10862), .C(n6419), .Y(
        \Decision_AXILiteS_s_axi_U/n834 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U752  ( .A(
        \Decision_AXILiteS_s_axi_U/n555 ), .B(n10863), .C(n6530), .Y(
        \Decision_AXILiteS_s_axi_U/n833 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U750  ( .A(
        \Decision_AXILiteS_s_axi_U/n555 ), .B(n10864), .C(n6642), .Y(
        \Decision_AXILiteS_s_axi_U/n832 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U748  ( .A(
        \Decision_AXILiteS_s_axi_U/n555 ), .B(n10865), .C(n6762), .Y(
        \Decision_AXILiteS_s_axi_U/n831 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U746  ( .A(
        \Decision_AXILiteS_s_axi_U/n555 ), .B(n10866), .C(n6889), .Y(
        \Decision_AXILiteS_s_axi_U/n830 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U744  ( .A(
        \Decision_AXILiteS_s_axi_U/n555 ), .B(n10867), .C(n7029), .Y(
        \Decision_AXILiteS_s_axi_U/n829 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U740  ( .A(n9305), .B(n7871), .C(n5032), 
        .Y(\Decision_AXILiteS_s_axi_U/n828 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U738  ( .A(n9304), .B(n7871), .C(n5031), 
        .Y(\Decision_AXILiteS_s_axi_U/n827 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U736  ( .A(n9303), .B(n7871), .C(n5030), 
        .Y(\Decision_AXILiteS_s_axi_U/n826 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U734  ( .A(n9302), .B(n7871), .C(n5029), 
        .Y(\Decision_AXILiteS_s_axi_U/n825 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U732  ( .A(n9301), .B(n7871), .C(n5028), 
        .Y(\Decision_AXILiteS_s_axi_U/n824 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U730  ( .A(n9300), .B(n7871), .C(n5027), 
        .Y(\Decision_AXILiteS_s_axi_U/n823 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U728  ( .A(n9299), .B(n7871), .C(n5026), 
        .Y(\Decision_AXILiteS_s_axi_U/n822 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U726  ( .A(n9298), .B(n7871), .C(n5025), 
        .Y(\Decision_AXILiteS_s_axi_U/n821 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U722  ( .A(n9297), .B(n8122), .C(n5024), 
        .Y(\Decision_AXILiteS_s_axi_U/n820 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U720  ( .A(n9296), .B(n8122), .C(n5023), 
        .Y(\Decision_AXILiteS_s_axi_U/n819 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U718  ( .A(n9295), .B(n8122), .C(n5022), 
        .Y(\Decision_AXILiteS_s_axi_U/n818 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U716  ( .A(n9294), .B(n8122), .C(n5021), 
        .Y(\Decision_AXILiteS_s_axi_U/n817 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U714  ( .A(n9293), .B(n8122), .C(n5020), 
        .Y(\Decision_AXILiteS_s_axi_U/n816 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U712  ( .A(n9292), .B(n8122), .C(n5019), 
        .Y(\Decision_AXILiteS_s_axi_U/n815 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U710  ( .A(n9291), .B(n8122), .C(n5018), 
        .Y(\Decision_AXILiteS_s_axi_U/n814 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U708  ( .A(n9290), .B(n8122), .C(n5017), 
        .Y(\Decision_AXILiteS_s_axi_U/n813 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U704  ( .A(n9289), .B(n8419), .C(n5016), 
        .Y(\Decision_AXILiteS_s_axi_U/n812 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U702  ( .A(n9288), .B(n8419), .C(n5015), 
        .Y(\Decision_AXILiteS_s_axi_U/n811 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U700  ( .A(n9287), .B(n8419), .C(n5014), 
        .Y(\Decision_AXILiteS_s_axi_U/n810 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U698  ( .A(n9286), .B(n8419), .C(n5013), 
        .Y(\Decision_AXILiteS_s_axi_U/n809 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U696  ( .A(n9285), .B(n8419), .C(n5012), 
        .Y(\Decision_AXILiteS_s_axi_U/n808 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U694  ( .A(n9284), .B(n8419), .C(n5011), 
        .Y(\Decision_AXILiteS_s_axi_U/n807 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U692  ( .A(n9283), .B(n8419), .C(n5010), 
        .Y(\Decision_AXILiteS_s_axi_U/n806 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U690  ( .A(n9282), .B(n8419), .C(n5009), 
        .Y(\Decision_AXILiteS_s_axi_U/n805 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U689  ( .A(n6810), .B(n5962), .C(ap_rst_n), .Y(\Decision_AXILiteS_s_axi_U/n492 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U687  ( .A(
        \Decision_AXILiteS_s_axi_U/n513 ), .B(n10852), .C(n6135), .Y(
        \Decision_AXILiteS_s_axi_U/n804 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U685  ( .A(
        \Decision_AXILiteS_s_axi_U/n513 ), .B(n10853), .C(n6216), .Y(
        \Decision_AXILiteS_s_axi_U/n803 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U683  ( .A(
        \Decision_AXILiteS_s_axi_U/n513 ), .B(n10854), .C(n6310), .Y(
        \Decision_AXILiteS_s_axi_U/n802 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U681  ( .A(
        \Decision_AXILiteS_s_axi_U/n513 ), .B(n10855), .C(n6418), .Y(
        \Decision_AXILiteS_s_axi_U/n801 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U679  ( .A(
        \Decision_AXILiteS_s_axi_U/n513 ), .B(n10856), .C(n6528), .Y(
        \Decision_AXILiteS_s_axi_U/n800 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U677  ( .A(
        \Decision_AXILiteS_s_axi_U/n513 ), .B(n10857), .C(n6640), .Y(
        \Decision_AXILiteS_s_axi_U/n799 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U675  ( .A(
        \Decision_AXILiteS_s_axi_U/n513 ), .B(n10858), .C(n7027), .Y(
        \Decision_AXILiteS_s_axi_U/n798 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U673  ( .A(
        \Decision_AXILiteS_s_axi_U/n513 ), .B(n10859), .C(n6887), .Y(
        \Decision_AXILiteS_s_axi_U/n797 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U669  ( .A(n9305), .B(n7656), .C(n5008), 
        .Y(\Decision_AXILiteS_s_axi_U/n796 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U667  ( .A(n9304), .B(n7656), .C(n5007), 
        .Y(\Decision_AXILiteS_s_axi_U/n795 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U665  ( .A(n9303), .B(n7656), .C(n5006), 
        .Y(\Decision_AXILiteS_s_axi_U/n794 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U663  ( .A(n9302), .B(n7656), .C(n5005), 
        .Y(\Decision_AXILiteS_s_axi_U/n793 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U661  ( .A(n9301), .B(n7656), .C(n5004), 
        .Y(\Decision_AXILiteS_s_axi_U/n792 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U659  ( .A(n9300), .B(n7656), .C(n5003), 
        .Y(\Decision_AXILiteS_s_axi_U/n791 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U657  ( .A(n9299), .B(n7656), .C(n5002), 
        .Y(\Decision_AXILiteS_s_axi_U/n790 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U655  ( .A(n9298), .B(n7656), .C(n5001), 
        .Y(\Decision_AXILiteS_s_axi_U/n789 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U651  ( .A(n9297), .B(n8418), .C(n5000), 
        .Y(\Decision_AXILiteS_s_axi_U/n788 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U649  ( .A(n9296), .B(n8418), .C(n4999), 
        .Y(\Decision_AXILiteS_s_axi_U/n787 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U647  ( .A(n9295), .B(n8418), .C(n4998), 
        .Y(\Decision_AXILiteS_s_axi_U/n786 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U645  ( .A(n9294), .B(n8418), .C(n4997), 
        .Y(\Decision_AXILiteS_s_axi_U/n785 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U643  ( .A(n9293), .B(n8418), .C(n4996), 
        .Y(\Decision_AXILiteS_s_axi_U/n784 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U641  ( .A(n9292), .B(n8418), .C(n4995), 
        .Y(\Decision_AXILiteS_s_axi_U/n783 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U639  ( .A(n9291), .B(n8418), .C(n4994), 
        .Y(\Decision_AXILiteS_s_axi_U/n782 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U637  ( .A(n9290), .B(n8418), .C(n4993), 
        .Y(\Decision_AXILiteS_s_axi_U/n781 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U633  ( .A(n9289), .B(n8121), .C(n6529), 
        .Y(\Decision_AXILiteS_s_axi_U/n780 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U631  ( .A(n9288), .B(n8121), .C(n6641), 
        .Y(\Decision_AXILiteS_s_axi_U/n779 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U629  ( .A(n9287), .B(n8121), .C(n6761), 
        .Y(\Decision_AXILiteS_s_axi_U/n778 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U627  ( .A(n9286), .B(n8121), .C(n6888), 
        .Y(\Decision_AXILiteS_s_axi_U/n777 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U625  ( .A(n9285), .B(n8121), .C(n7028), 
        .Y(\Decision_AXILiteS_s_axi_U/n776 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U623  ( .A(n9284), .B(n8121), .C(n7182), 
        .Y(\Decision_AXILiteS_s_axi_U/n775 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U621  ( .A(n9283), .B(n8121), .C(n7345), 
        .Y(\Decision_AXILiteS_s_axi_U/n774 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U619  ( .A(n9282), .B(n8121), .C(n7524), 
        .Y(\Decision_AXILiteS_s_axi_U/n773 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U618  ( .A(
        \Decision_AXILiteS_s_axi_U/n371 ), .B(n10898), .C(
        \Decision_AXILiteS_s_axi_U/waddr[6] ), .Y(
        \Decision_AXILiteS_s_axi_U/n418 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U617  ( .A(n7258), .B(n7434), .C(ap_rst_n), .Y(\Decision_AXILiteS_s_axi_U/n473 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U615  ( .A(
        \Decision_AXILiteS_s_axi_U/n471 ), .B(n10844), .C(n4992), .Y(
        \Decision_AXILiteS_s_axi_U/n772 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U613  ( .A(
        \Decision_AXILiteS_s_axi_U/n471 ), .B(n10845), .C(n4991), .Y(
        \Decision_AXILiteS_s_axi_U/n771 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U611  ( .A(
        \Decision_AXILiteS_s_axi_U/n471 ), .B(n10846), .C(n4990), .Y(
        \Decision_AXILiteS_s_axi_U/n770 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U609  ( .A(
        \Decision_AXILiteS_s_axi_U/n471 ), .B(n10847), .C(n4989), .Y(
        \Decision_AXILiteS_s_axi_U/n769 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U607  ( .A(
        \Decision_AXILiteS_s_axi_U/n471 ), .B(n10848), .C(n4988), .Y(
        \Decision_AXILiteS_s_axi_U/n768 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U605  ( .A(
        \Decision_AXILiteS_s_axi_U/n471 ), .B(n10849), .C(n4987), .Y(
        \Decision_AXILiteS_s_axi_U/n767 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U603  ( .A(
        \Decision_AXILiteS_s_axi_U/n471 ), .B(n10850), .C(n4986), .Y(
        \Decision_AXILiteS_s_axi_U/n766 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U601  ( .A(
        \Decision_AXILiteS_s_axi_U/n471 ), .B(n10851), .C(n4985), .Y(
        \Decision_AXILiteS_s_axi_U/n765 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U600  ( .A(
        \Decision_AXILiteS_s_axi_U/waddr[3] ), .B(n10897), .C(n9279), .Y(
        \Decision_AXILiteS_s_axi_U/n470 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U597  ( .A(
        \Decision_AXILiteS_s_axi_U/n460 ), .B(n10836), .C(n6760), .Y(
        \Decision_AXILiteS_s_axi_U/n764 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U595  ( .A(
        \Decision_AXILiteS_s_axi_U/n460 ), .B(n10837), .C(n6886), .Y(
        \Decision_AXILiteS_s_axi_U/n763 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U593  ( .A(
        \Decision_AXILiteS_s_axi_U/n460 ), .B(n10838), .C(n7026), .Y(
        \Decision_AXILiteS_s_axi_U/n762 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U591  ( .A(
        \Decision_AXILiteS_s_axi_U/n460 ), .B(n10839), .C(n7181), .Y(
        \Decision_AXILiteS_s_axi_U/n761 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U589  ( .A(
        \Decision_AXILiteS_s_axi_U/n460 ), .B(n10840), .C(n7344), .Y(
        \Decision_AXILiteS_s_axi_U/n760 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U587  ( .A(
        \Decision_AXILiteS_s_axi_U/n460 ), .B(n10841), .C(n7523), .Y(
        \Decision_AXILiteS_s_axi_U/n759 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U585  ( .A(
        \Decision_AXILiteS_s_axi_U/n460 ), .B(n10842), .C(n7722), .Y(
        \Decision_AXILiteS_s_axi_U/n758 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U583  ( .A(
        \Decision_AXILiteS_s_axi_U/n460 ), .B(n10843), .C(n7939), .Y(
        \Decision_AXILiteS_s_axi_U/n757 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U582  ( .A(
        \Decision_AXILiteS_s_axi_U/waddr[4] ), .B(n10895), .C(n9279), .Y(
        \Decision_AXILiteS_s_axi_U/n459 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U579  ( .A(
        \Decision_AXILiteS_s_axi_U/n450 ), .B(n10828), .C(n6309), .Y(
        \Decision_AXILiteS_s_axi_U/n756 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U577  ( .A(
        \Decision_AXILiteS_s_axi_U/n450 ), .B(n10829), .C(n6416), .Y(
        \Decision_AXILiteS_s_axi_U/n755 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U575  ( .A(
        \Decision_AXILiteS_s_axi_U/n450 ), .B(n10830), .C(n6215), .Y(
        \Decision_AXILiteS_s_axi_U/n754 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U573  ( .A(
        \Decision_AXILiteS_s_axi_U/n450 ), .B(n10831), .C(n6639), .Y(
        \Decision_AXILiteS_s_axi_U/n753 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U571  ( .A(
        \Decision_AXILiteS_s_axi_U/n450 ), .B(n10832), .C(n6758), .Y(
        \Decision_AXILiteS_s_axi_U/n752 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U569  ( .A(
        \Decision_AXILiteS_s_axi_U/n450 ), .B(n10833), .C(n6526), .Y(
        \Decision_AXILiteS_s_axi_U/n751 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U567  ( .A(
        \Decision_AXILiteS_s_axi_U/n450 ), .B(n10834), .C(n7179), .Y(
        \Decision_AXILiteS_s_axi_U/n750 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U565  ( .A(
        \Decision_AXILiteS_s_axi_U/n450 ), .B(n10835), .C(n7342), .Y(
        \Decision_AXILiteS_s_axi_U/n749 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U561  ( .A(n9305), .B(n8417), .C(n4984), 
        .Y(\Decision_AXILiteS_s_axi_U/n748 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U559  ( .A(n9304), .B(n8417), .C(n4983), 
        .Y(\Decision_AXILiteS_s_axi_U/n747 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U557  ( .A(n9303), .B(n8417), .C(n4982), 
        .Y(\Decision_AXILiteS_s_axi_U/n746 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U555  ( .A(n9302), .B(n8417), .C(n4981), 
        .Y(\Decision_AXILiteS_s_axi_U/n745 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U553  ( .A(n9301), .B(n8417), .C(n4980), 
        .Y(\Decision_AXILiteS_s_axi_U/n744 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U551  ( .A(n9300), .B(n8417), .C(n4979), 
        .Y(\Decision_AXILiteS_s_axi_U/n743 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U549  ( .A(n9299), .B(n8417), .C(n4978), 
        .Y(\Decision_AXILiteS_s_axi_U/n742 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U547  ( .A(n9298), .B(n8417), .C(n4977), 
        .Y(\Decision_AXILiteS_s_axi_U/n741 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U543  ( .A(n9297), .B(n7655), .C(n4976), 
        .Y(\Decision_AXILiteS_s_axi_U/n740 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U541  ( .A(n9296), .B(n7655), .C(n4975), 
        .Y(\Decision_AXILiteS_s_axi_U/n739 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U539  ( .A(n9295), .B(n7655), .C(n4974), 
        .Y(\Decision_AXILiteS_s_axi_U/n738 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U537  ( .A(n9294), .B(n7655), .C(n4973), 
        .Y(\Decision_AXILiteS_s_axi_U/n737 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U535  ( .A(n9293), .B(n7655), .C(n4972), 
        .Y(\Decision_AXILiteS_s_axi_U/n736 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U533  ( .A(n9292), .B(n7655), .C(n4971), 
        .Y(\Decision_AXILiteS_s_axi_U/n735 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U531  ( .A(n9291), .B(n7655), .C(n4970), 
        .Y(\Decision_AXILiteS_s_axi_U/n734 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U529  ( .A(n9290), .B(n7655), .C(n4969), 
        .Y(\Decision_AXILiteS_s_axi_U/n733 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U525  ( .A(n9289), .B(n7870), .C(n6417), 
        .Y(\Decision_AXILiteS_s_axi_U/n732 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U523  ( .A(n9288), .B(n7870), .C(n6527), 
        .Y(\Decision_AXILiteS_s_axi_U/n731 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U521  ( .A(n9287), .B(n7870), .C(n6885), 
        .Y(\Decision_AXILiteS_s_axi_U/n730 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U519  ( .A(n9286), .B(n7870), .C(n6759), 
        .Y(\Decision_AXILiteS_s_axi_U/n729 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U517  ( .A(n9285), .B(n7870), .C(n7180), 
        .Y(\Decision_AXILiteS_s_axi_U/n728 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U515  ( .A(n9284), .B(n7870), .C(n7025), 
        .Y(\Decision_AXILiteS_s_axi_U/n727 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U513  ( .A(n9283), .B(n7870), .C(n7522), 
        .Y(\Decision_AXILiteS_s_axi_U/n726 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U511  ( .A(n9282), .B(n7870), .C(n7343), 
        .Y(\Decision_AXILiteS_s_axi_U/n725 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U510  ( .A(n6810), .B(n7434), .C(ap_rst_n), .Y(\Decision_AXILiteS_s_axi_U/n383 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U508  ( .A(
        \Decision_AXILiteS_s_axi_U/n408 ), .B(n10820), .C(n6068), .Y(
        \Decision_AXILiteS_s_axi_U/n724 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U506  ( .A(
        \Decision_AXILiteS_s_axi_U/n408 ), .B(n10821), .C(n6134), .Y(
        \Decision_AXILiteS_s_axi_U/n723 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U504  ( .A(
        \Decision_AXILiteS_s_axi_U/n408 ), .B(n10822), .C(n6525), .Y(
        \Decision_AXILiteS_s_axi_U/n722 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U502  ( .A(
        \Decision_AXILiteS_s_axi_U/n408 ), .B(n10823), .C(n6214), .Y(
        \Decision_AXILiteS_s_axi_U/n721 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U500  ( .A(
        \Decision_AXILiteS_s_axi_U/n408 ), .B(n10824), .C(n6308), .Y(
        \Decision_AXILiteS_s_axi_U/n720 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U498  ( .A(
        \Decision_AXILiteS_s_axi_U/n408 ), .B(n10825), .C(n6415), .Y(
        \Decision_AXILiteS_s_axi_U/n719 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U496  ( .A(
        \Decision_AXILiteS_s_axi_U/n408 ), .B(n10826), .C(n6638), .Y(
        \Decision_AXILiteS_s_axi_U/n718 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U494  ( .A(
        \Decision_AXILiteS_s_axi_U/n408 ), .B(n10827), .C(n7177), .Y(
        \Decision_AXILiteS_s_axi_U/n717 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U490  ( .A(n9305), .B(n8120), .C(n4968), 
        .Y(\Decision_AXILiteS_s_axi_U/n716 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U488  ( .A(n9304), .B(n8120), .C(n4967), 
        .Y(\Decision_AXILiteS_s_axi_U/n715 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U486  ( .A(n9303), .B(n8120), .C(n4966), 
        .Y(\Decision_AXILiteS_s_axi_U/n714 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U484  ( .A(n9302), .B(n8120), .C(n4965), 
        .Y(\Decision_AXILiteS_s_axi_U/n713 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U482  ( .A(n9301), .B(n8120), .C(n4964), 
        .Y(\Decision_AXILiteS_s_axi_U/n712 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U480  ( .A(n9300), .B(n8120), .C(n4963), 
        .Y(\Decision_AXILiteS_s_axi_U/n711 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U478  ( .A(n9299), .B(n8120), .C(n4962), 
        .Y(\Decision_AXILiteS_s_axi_U/n710 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U476  ( .A(n9298), .B(n8120), .C(n4961), 
        .Y(\Decision_AXILiteS_s_axi_U/n709 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U472  ( .A(n7866), .B(n9297), .C(n4960), 
        .Y(\Decision_AXILiteS_s_axi_U/n708 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U470  ( .A(n7866), .B(n9296), .C(n4959), 
        .Y(\Decision_AXILiteS_s_axi_U/n707 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U468  ( .A(n7866), .B(n9295), .C(n4958), 
        .Y(\Decision_AXILiteS_s_axi_U/n706 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U466  ( .A(n7866), .B(n9294), .C(n4957), 
        .Y(\Decision_AXILiteS_s_axi_U/n705 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U464  ( .A(n7866), .B(n9293), .C(n4956), 
        .Y(\Decision_AXILiteS_s_axi_U/n704 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U462  ( .A(n7866), .B(n9292), .C(n4955), 
        .Y(\Decision_AXILiteS_s_axi_U/n703 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U460  ( .A(n7866), .B(n9291), .C(n4954), 
        .Y(\Decision_AXILiteS_s_axi_U/n702 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U458  ( .A(n7866), .B(n9290), .C(n4953), 
        .Y(\Decision_AXILiteS_s_axi_U/n701 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U454  ( .A(n7652), .B(n9289), .C(n4952), 
        .Y(\Decision_AXILiteS_s_axi_U/n700 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U452  ( .A(n7652), .B(n9288), .C(n4951), 
        .Y(\Decision_AXILiteS_s_axi_U/n699 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U450  ( .A(n7652), .B(n9287), .C(n4950), 
        .Y(\Decision_AXILiteS_s_axi_U/n698 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U448  ( .A(n7652), .B(n9286), .C(n4949), 
        .Y(\Decision_AXILiteS_s_axi_U/n697 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U446  ( .A(n7652), .B(n9285), .C(n4948), 
        .Y(\Decision_AXILiteS_s_axi_U/n696 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U444  ( .A(n7652), .B(n9284), .C(n7341), 
        .Y(\Decision_AXILiteS_s_axi_U/n695 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U442  ( .A(n7652), .B(n9283), .C(n4947), 
        .Y(\Decision_AXILiteS_s_axi_U/n694 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U440  ( .A(n7652), .B(n9282), .C(n7178), 
        .Y(\Decision_AXILiteS_s_axi_U/n693 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U438  ( .A(
        \Decision_AXILiteS_s_axi_U/n371 ), .B(\Decision_AXILiteS_s_axi_U/n481 ), .C(n7084), .Y(\Decision_AXILiteS_s_axi_U/n370 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U435  ( .A(
        \Decision_AXILiteS_s_axi_U/n354 ), .B(n10812), .C(n6524), .Y(
        \Decision_AXILiteS_s_axi_U/n692 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U433  ( .A(
        \Decision_AXILiteS_s_axi_U/n354 ), .B(n10813), .C(n6637), .Y(
        \Decision_AXILiteS_s_axi_U/n691 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U431  ( .A(
        \Decision_AXILiteS_s_axi_U/n354 ), .B(n10814), .C(n6757), .Y(
        \Decision_AXILiteS_s_axi_U/n690 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U429  ( .A(
        \Decision_AXILiteS_s_axi_U/n354 ), .B(n10815), .C(n6884), .Y(
        \Decision_AXILiteS_s_axi_U/n689 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U427  ( .A(
        \Decision_AXILiteS_s_axi_U/n354 ), .B(n10816), .C(n7521), .Y(
        \Decision_AXILiteS_s_axi_U/n688 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U425  ( .A(
        \Decision_AXILiteS_s_axi_U/n354 ), .B(n10817), .C(n7176), .Y(
        \Decision_AXILiteS_s_axi_U/n687 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U423  ( .A(
        \Decision_AXILiteS_s_axi_U/n354 ), .B(n10818), .C(n7938), .Y(
        \Decision_AXILiteS_s_axi_U/n686 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U421  ( .A(
        \Decision_AXILiteS_s_axi_U/n354 ), .B(n10819), .C(n7721), .Y(
        \Decision_AXILiteS_s_axi_U/n685 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U417  ( .A(n7447), .B(n9305), .C(n4946), 
        .Y(\Decision_AXILiteS_s_axi_U/n684 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U415  ( .A(n7447), .B(n9304), .C(n4945), 
        .Y(\Decision_AXILiteS_s_axi_U/n683 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U413  ( .A(n7447), .B(n9303), .C(n4944), 
        .Y(\Decision_AXILiteS_s_axi_U/n682 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U411  ( .A(n7447), .B(n9302), .C(n4943), 
        .Y(\Decision_AXILiteS_s_axi_U/n681 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U409  ( .A(n7447), .B(n9301), .C(n4942), 
        .Y(\Decision_AXILiteS_s_axi_U/n680 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U407  ( .A(n7447), .B(n9300), .C(n4941), 
        .Y(\Decision_AXILiteS_s_axi_U/n679 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U405  ( .A(n7447), .B(n9299), .C(n4940), 
        .Y(\Decision_AXILiteS_s_axi_U/n678 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U403  ( .A(n7447), .B(n9298), .C(n4939), 
        .Y(\Decision_AXILiteS_s_axi_U/n677 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U400  ( .A(n9321), .B(n9317), .C(
        s_axi_AXILiteS_ARADDR[4]), .Y(\Decision_AXILiteS_s_axi_U/n319 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U399  ( .A(n9311), .B(n9320), .C(n8859), 
        .Y(\Decision_AXILiteS_s_axi_U/n340 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U398  ( .A(n8859), .B(n9311), .C(n8858), 
        .Y(\Decision_AXILiteS_s_axi_U/n339 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U397  ( .A(athresh[0]), .B(n9309), .C(
        vthresh[0]), .D(n9310), .Y(\Decision_AXILiteS_s_axi_U/n326 ) );
  NOR3X1 \Decision_AXILiteS_s_axi_U/U396  ( .A(n8857), .B(n8859), .C(n9317), 
        .Y(\Decision_AXILiteS_s_axi_U/n321 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U395  ( .A(s_axi_AXILiteS_ARADDR[4]), .B(
        n9320), .C(\Decision_AXILiteS_s_axi_U/n321 ), .Y(
        \Decision_AXILiteS_s_axi_U/n338 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U392  ( .A(
        \Decision_AXILiteS_s_axi_U/int_ier[0] ), .B(n9321), .C(
        \Decision_AXILiteS_s_axi_U/int_isr[0] ), .D(n8857), .Y(
        \Decision_AXILiteS_s_axi_U/n336 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U391  ( .A(n8857), .B(n9320), .C(
        \Decision_AXILiteS_s_axi_U/int_gie ), .Y(
        \Decision_AXILiteS_s_axi_U/n337 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U390  ( .A(n5531), .B(n9320), .C(n4920), 
        .Y(\Decision_AXILiteS_s_axi_U/n335 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U389  ( .A(n7999), .B(\reset_A_V[0] ), 
        .C(\Decision_AXILiteS_s_axi_U/n310 ), .D(
        \Decision_AXILiteS_s_axi_U/n335 ), .Y(\Decision_AXILiteS_s_axi_U/n330 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U388  ( .A(\reset_V_V[0] ), .B(n9320), 
        .C(\reset_params_V[0] ), .D(n8858), .Y(
        \Decision_AXILiteS_s_axi_U/n333 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U386  ( .A(
        \Decision_AXILiteS_s_axi_U/n310 ), .B(n8859), .C(n8267), .Y(
        \Decision_AXILiteS_s_axi_U/n331 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U385  ( .A(n8859), .B(n5699), .C(n4919), 
        .Y(\Decision_AXILiteS_s_axi_U/n329 ) );
  AOI21X1 \Decision_AXILiteS_s_axi_U/U384  ( .A(ap_start), .B(n9316), .C(
        \Decision_AXILiteS_s_axi_U/n329 ), .Y(\Decision_AXILiteS_s_axi_U/n328 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U383  ( .A(n5449), .B(n5693), .C(n5875), 
        .Y(\Decision_AXILiteS_s_axi_U/n313 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U382  ( .A(n8858), .B(
        s_axi_AXILiteS_ARADDR[4]), .C(\Decision_AXILiteS_s_axi_U/n321 ), .Y(
        \Decision_AXILiteS_s_axi_U/n325 ) );
  NOR3X1 \Decision_AXILiteS_s_axi_U/U381  ( .A(n8857), .B(
        s_axi_AXILiteS_ARADDR[4]), .C(n8858), .Y(
        \Decision_AXILiteS_s_axi_U/n324 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U380  ( .A(s_axi_AXILiteS_ARADDR[6]), .B(
        n8859), .C(\Decision_AXILiteS_s_axi_U/n324 ), .Y(
        \Decision_AXILiteS_s_axi_U/n323 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U379  ( .A(v_length[0]), .B(n9313), .C(
        data[0]), .D(n9318), .Y(\Decision_AXILiteS_s_axi_U/n316 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U378  ( .A(n8858), .B(n9319), .C(
        \Decision_AXILiteS_s_axi_U/n321 ), .Y(\Decision_AXILiteS_s_axi_U/n322 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U376  ( .A(n9320), .B(n9319), .C(
        \Decision_AXILiteS_s_axi_U/n321 ), .Y(\Decision_AXILiteS_s_axi_U/n320 ) );
  NOR3X1 \Decision_AXILiteS_s_axi_U/U375  ( .A(n8858), .B(n8859), .C(n8383), 
        .Y(\Decision_AXILiteS_s_axi_U/n247 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U374  ( .A(a_flip[0]), .B(n9315), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[0] ), .D(
        \Decision_AXILiteS_s_axi_U/n247 ), .Y(\Decision_AXILiteS_s_axi_U/n318 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U371  ( .A(n5547), .B(n5715), .C(
        \Decision_AXILiteS_s_axi_U/n248 ), .Y(\Decision_AXILiteS_s_axi_U/n312 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U367  ( .A(
        \Decision_AXILiteS_s_axi_U/int_ier[1] ), .B(n9321), .C(
        \Decision_AXILiteS_s_axi_U/int_isr[1] ), .D(n8857), .Y(
        \Decision_AXILiteS_s_axi_U/n309 ) );
  NOR3X1 \Decision_AXILiteS_s_axi_U/U366  ( .A(n5898), .B(n8859), .C(n5904), 
        .Y(\Decision_AXILiteS_s_axi_U/n307 ) );
  AOI21X1 \Decision_AXILiteS_s_axi_U/U365  ( .A(
        \Decision_AXILiteS_s_axi_U/int_ap_done ), .B(n9316), .C(
        \Decision_AXILiteS_s_axi_U/n307 ), .Y(\Decision_AXILiteS_s_axi_U/n304 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U363  ( .A(vthresh[1]), .B(n9310), .C(
        a_length[1]), .D(n9312), .Y(\Decision_AXILiteS_s_axi_U/n306 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U362  ( .A(n5482), .B(n5692), .C(n5856), 
        .Y(\Decision_AXILiteS_s_axi_U/n299 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U361  ( .A(v_length[1]), .B(n9313), .C(
        data[1]), .D(n9318), .Y(\Decision_AXILiteS_s_axi_U/n301 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U359  ( .A(a_flip[1]), .B(n9315), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[1] ), .D(
        \Decision_AXILiteS_s_axi_U/n247 ), .Y(\Decision_AXILiteS_s_axi_U/n303 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U357  ( .A(n5546), .B(n5712), .C(
        \Decision_AXILiteS_s_axi_U/n248 ), .Y(\Decision_AXILiteS_s_axi_U/n298 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U354  ( .A(n2154), .B(n9316), .C(
        athresh[2]), .D(n9309), .Y(\Decision_AXILiteS_s_axi_U/n294 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U352  ( .A(a_length[2]), .B(n9312), .C(
        v_length[2]), .D(n9313), .Y(\Decision_AXILiteS_s_axi_U/n296 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U351  ( .A(n5448), .B(n5691), .C(n5853), 
        .Y(\Decision_AXILiteS_s_axi_U/n290 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U350  ( .A(a_flip[2]), .B(n9315), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[2] ), .D(
        \Decision_AXILiteS_s_axi_U/n247 ), .Y(\Decision_AXILiteS_s_axi_U/n292 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U349  ( .A(data[2]), .B(n9318), .C(
        v_flip[2]), .D(n9314), .Y(\Decision_AXILiteS_s_axi_U/n293 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U347  ( .A(n5545), .B(n5721), .C(
        \Decision_AXILiteS_s_axi_U/n248 ), .Y(\Decision_AXILiteS_s_axi_U/n289 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U344  ( .A(n9316), .B(ap_CS_fsm[13]), .C(
        athresh[3]), .D(n9309), .Y(\Decision_AXILiteS_s_axi_U/n285 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U342  ( .A(a_length[3]), .B(n9312), .C(
        v_length[3]), .D(n9313), .Y(\Decision_AXILiteS_s_axi_U/n287 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U341  ( .A(n5447), .B(n5690), .C(n5852), 
        .Y(\Decision_AXILiteS_s_axi_U/n281 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U340  ( .A(a_flip[3]), .B(n9315), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[3] ), .D(
        \Decision_AXILiteS_s_axi_U/n247 ), .Y(\Decision_AXILiteS_s_axi_U/n283 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U339  ( .A(data[3]), .B(n9318), .C(
        v_flip[3]), .D(n9314), .Y(\Decision_AXILiteS_s_axi_U/n284 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U337  ( .A(n5544), .B(n5720), .C(
        \Decision_AXILiteS_s_axi_U/n248 ), .Y(\Decision_AXILiteS_s_axi_U/n280 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U335  ( .A(a_flip[4]), .B(n9315), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[4] ), .D(
        \Decision_AXILiteS_s_axi_U/n247 ), .Y(\Decision_AXILiteS_s_axi_U/n274 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U334  ( .A(data[4]), .B(n9318), .C(
        v_flip[4]), .D(n9314), .Y(\Decision_AXILiteS_s_axi_U/n275 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U333  ( .A(a_length[4]), .B(n9312), .C(
        v_length[4]), .D(n9313), .Y(\Decision_AXILiteS_s_axi_U/n277 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U332  ( .A(athresh[4]), .B(n9309), .C(
        vthresh[4]), .D(n9310), .Y(\Decision_AXILiteS_s_axi_U/n278 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U331  ( .A(n5446), .B(n5566), .C(
        \Decision_AXILiteS_s_axi_U/n276 ), .Y(\Decision_AXILiteS_s_axi_U/n273 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U330  ( .A(
        \Decision_AXILiteS_s_axi_U/n248 ), .B(n5561), .C(
        s_axi_AXILiteS_RDATA[4]), .D(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n272 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U329  ( .A(a_flip[5]), .B(n9315), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[5] ), .D(
        \Decision_AXILiteS_s_axi_U/n247 ), .Y(\Decision_AXILiteS_s_axi_U/n267 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U328  ( .A(data[5]), .B(n9318), .C(
        v_flip[5]), .D(n9314), .Y(\Decision_AXILiteS_s_axi_U/n268 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U327  ( .A(a_length[5]), .B(n9312), .C(
        v_length[5]), .D(n9313), .Y(\Decision_AXILiteS_s_axi_U/n270 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U326  ( .A(athresh[5]), .B(n9309), .C(
        vthresh[5]), .D(n9310), .Y(\Decision_AXILiteS_s_axi_U/n271 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U325  ( .A(n5445), .B(n5565), .C(
        \Decision_AXILiteS_s_axi_U/n269 ), .Y(\Decision_AXILiteS_s_axi_U/n266 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U324  ( .A(
        \Decision_AXILiteS_s_axi_U/n248 ), .B(n5560), .C(
        s_axi_AXILiteS_RDATA[5]), .D(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n265 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U323  ( .A(a_flip[6]), .B(n9315), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[6] ), .D(
        \Decision_AXILiteS_s_axi_U/n247 ), .Y(\Decision_AXILiteS_s_axi_U/n260 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U322  ( .A(data[6]), .B(n9318), .C(
        v_flip[6]), .D(n9314), .Y(\Decision_AXILiteS_s_axi_U/n261 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U321  ( .A(a_length[6]), .B(n9312), .C(
        v_length[6]), .D(n9313), .Y(\Decision_AXILiteS_s_axi_U/n263 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U320  ( .A(athresh[6]), .B(n9309), .C(
        vthresh[6]), .D(n9310), .Y(\Decision_AXILiteS_s_axi_U/n264 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U319  ( .A(n5444), .B(n5564), .C(
        \Decision_AXILiteS_s_axi_U/n262 ), .Y(\Decision_AXILiteS_s_axi_U/n259 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U318  ( .A(
        \Decision_AXILiteS_s_axi_U/n248 ), .B(n5559), .C(
        s_axi_AXILiteS_RDATA[6]), .D(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n258 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U316  ( .A(
        \Decision_AXILiteS_s_axi_U/int_auto_restart ), .B(n9316), .C(
        athresh[7]), .D(n9309), .Y(\Decision_AXILiteS_s_axi_U/n255 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U314  ( .A(a_length[7]), .B(n9312), .C(
        v_length[7]), .D(n9313), .Y(\Decision_AXILiteS_s_axi_U/n257 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U313  ( .A(n5443), .B(n5689), .C(n5851), 
        .Y(\Decision_AXILiteS_s_axi_U/n251 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U312  ( .A(a_flip[7]), .B(n9315), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[7] ), .D(
        \Decision_AXILiteS_s_axi_U/n247 ), .Y(\Decision_AXILiteS_s_axi_U/n253 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U311  ( .A(data[7]), .B(n9318), .C(
        v_flip[7]), .D(n9314), .Y(\Decision_AXILiteS_s_axi_U/n254 ) );
  OAI21X1 \Decision_AXILiteS_s_axi_U/U309  ( .A(n5543), .B(n5719), .C(
        \Decision_AXILiteS_s_axi_U/n248 ), .Y(\Decision_AXILiteS_s_axi_U/n250 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U307  ( .A(a_length[8]), .B(
        \Decision_AXILiteS_s_axi_U/n157 ), .C(v_length[8]), .D(
        \Decision_AXILiteS_s_axi_U/n155 ), .Y(\Decision_AXILiteS_s_axi_U/n242 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U305  ( .A(athresh[8]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[8]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n245 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U304  ( .A(data[8]), .B(
        \Decision_AXILiteS_s_axi_U/n210 ), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[8] ), .D(
        \Decision_AXILiteS_s_axi_U/n211 ), .Y(\Decision_AXILiteS_s_axi_U/n246 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U303  ( .A(n5442), .B(n5688), .C(
        \Decision_AXILiteS_s_axi_U/n244 ), .Y(\Decision_AXILiteS_s_axi_U/n671 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U302  ( .A(a_length[9]), .B(
        \Decision_AXILiteS_s_axi_U/n157 ), .C(v_length[9]), .D(
        \Decision_AXILiteS_s_axi_U/n155 ), .Y(\Decision_AXILiteS_s_axi_U/n237 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U300  ( .A(athresh[9]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[9]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n240 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U299  ( .A(data[9]), .B(
        \Decision_AXILiteS_s_axi_U/n210 ), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[9] ), .D(
        \Decision_AXILiteS_s_axi_U/n211 ), .Y(\Decision_AXILiteS_s_axi_U/n241 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U298  ( .A(n5441), .B(n5687), .C(
        \Decision_AXILiteS_s_axi_U/n239 ), .Y(\Decision_AXILiteS_s_axi_U/n670 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U297  ( .A(a_length[10]), .B(
        \Decision_AXILiteS_s_axi_U/n157 ), .C(v_length[10]), .D(
        \Decision_AXILiteS_s_axi_U/n155 ), .Y(\Decision_AXILiteS_s_axi_U/n232 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U295  ( .A(athresh[10]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[10]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n235 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U294  ( .A(data[10]), .B(
        \Decision_AXILiteS_s_axi_U/n210 ), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[10] ), .D(
        \Decision_AXILiteS_s_axi_U/n211 ), .Y(\Decision_AXILiteS_s_axi_U/n236 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U293  ( .A(n5440), .B(n5686), .C(
        \Decision_AXILiteS_s_axi_U/n234 ), .Y(\Decision_AXILiteS_s_axi_U/n669 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U292  ( .A(a_length[11]), .B(
        \Decision_AXILiteS_s_axi_U/n157 ), .C(v_length[11]), .D(
        \Decision_AXILiteS_s_axi_U/n155 ), .Y(\Decision_AXILiteS_s_axi_U/n227 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U290  ( .A(athresh[11]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[11]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n230 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U289  ( .A(data[11]), .B(
        \Decision_AXILiteS_s_axi_U/n210 ), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[11] ), .D(
        \Decision_AXILiteS_s_axi_U/n211 ), .Y(\Decision_AXILiteS_s_axi_U/n231 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U288  ( .A(n5439), .B(n5685), .C(
        \Decision_AXILiteS_s_axi_U/n229 ), .Y(\Decision_AXILiteS_s_axi_U/n668 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U287  ( .A(a_length[12]), .B(
        \Decision_AXILiteS_s_axi_U/n157 ), .C(v_length[12]), .D(
        \Decision_AXILiteS_s_axi_U/n155 ), .Y(\Decision_AXILiteS_s_axi_U/n222 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U285  ( .A(athresh[12]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[12]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n225 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U284  ( .A(data[12]), .B(
        \Decision_AXILiteS_s_axi_U/n210 ), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[12] ), .D(
        \Decision_AXILiteS_s_axi_U/n211 ), .Y(\Decision_AXILiteS_s_axi_U/n226 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U283  ( .A(n5438), .B(n5684), .C(
        \Decision_AXILiteS_s_axi_U/n224 ), .Y(\Decision_AXILiteS_s_axi_U/n667 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U282  ( .A(a_length[13]), .B(
        \Decision_AXILiteS_s_axi_U/n157 ), .C(v_length[13]), .D(
        \Decision_AXILiteS_s_axi_U/n155 ), .Y(\Decision_AXILiteS_s_axi_U/n217 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U280  ( .A(athresh[13]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[13]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n220 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U279  ( .A(data[13]), .B(
        \Decision_AXILiteS_s_axi_U/n210 ), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[13] ), .D(
        \Decision_AXILiteS_s_axi_U/n211 ), .Y(\Decision_AXILiteS_s_axi_U/n221 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U278  ( .A(n5437), .B(n5683), .C(
        \Decision_AXILiteS_s_axi_U/n219 ), .Y(\Decision_AXILiteS_s_axi_U/n666 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U277  ( .A(a_length[14]), .B(
        \Decision_AXILiteS_s_axi_U/n157 ), .C(v_length[14]), .D(
        \Decision_AXILiteS_s_axi_U/n155 ), .Y(\Decision_AXILiteS_s_axi_U/n212 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U275  ( .A(athresh[14]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[14]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n215 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U274  ( .A(data[14]), .B(
        \Decision_AXILiteS_s_axi_U/n210 ), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[14] ), .D(
        \Decision_AXILiteS_s_axi_U/n211 ), .Y(\Decision_AXILiteS_s_axi_U/n216 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U273  ( .A(n5436), .B(n5682), .C(
        \Decision_AXILiteS_s_axi_U/n214 ), .Y(\Decision_AXILiteS_s_axi_U/n665 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U272  ( .A(a_length[15]), .B(
        \Decision_AXILiteS_s_axi_U/n157 ), .C(v_length[15]), .D(
        \Decision_AXILiteS_s_axi_U/n155 ), .Y(\Decision_AXILiteS_s_axi_U/n205 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U270  ( .A(athresh[15]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[15]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n208 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U269  ( .A(data[15]), .B(
        \Decision_AXILiteS_s_axi_U/n210 ), .C(
        \Decision_AXILiteS_s_axi_U/int_ap_return[15] ), .D(
        \Decision_AXILiteS_s_axi_U/n211 ), .Y(\Decision_AXILiteS_s_axi_U/n209 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U268  ( .A(n5435), .B(n5681), .C(
        \Decision_AXILiteS_s_axi_U/n207 ), .Y(\Decision_AXILiteS_s_axi_U/n664 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U267  ( .A(athresh[16]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[16]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n202 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U265  ( .A(v_length[16]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[16]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n204 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U264  ( .A(n5434), .B(n5680), .C(n5850), 
        .Y(\Decision_AXILiteS_s_axi_U/n663 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U263  ( .A(athresh[17]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[17]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n199 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U261  ( .A(v_length[17]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[17]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n201 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U260  ( .A(n5433), .B(n5679), .C(n5849), 
        .Y(\Decision_AXILiteS_s_axi_U/n662 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U259  ( .A(athresh[18]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[18]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n196 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U257  ( .A(v_length[18]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[18]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n198 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U256  ( .A(n5432), .B(n5678), .C(n5848), 
        .Y(\Decision_AXILiteS_s_axi_U/n661 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U255  ( .A(athresh[19]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[19]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n193 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U253  ( .A(v_length[19]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[19]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n195 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U252  ( .A(n5431), .B(n5677), .C(n5847), 
        .Y(\Decision_AXILiteS_s_axi_U/n660 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U251  ( .A(athresh[20]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[20]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n190 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U249  ( .A(v_length[20]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[20]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n192 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U248  ( .A(n5430), .B(n5676), .C(n5846), 
        .Y(\Decision_AXILiteS_s_axi_U/n659 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U247  ( .A(athresh[21]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[21]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n187 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U245  ( .A(v_length[21]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[21]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n189 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U244  ( .A(n5429), .B(n5675), .C(n5845), 
        .Y(\Decision_AXILiteS_s_axi_U/n658 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U243  ( .A(athresh[22]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[22]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n184 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U241  ( .A(v_length[22]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[22]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n186 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U240  ( .A(n5428), .B(n5674), .C(n5844), 
        .Y(\Decision_AXILiteS_s_axi_U/n657 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U239  ( .A(athresh[23]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[23]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n181 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U237  ( .A(v_length[23]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[23]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n183 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U236  ( .A(n5427), .B(n5673), .C(n5843), 
        .Y(\Decision_AXILiteS_s_axi_U/n656 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U235  ( .A(athresh[24]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[24]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n178 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U233  ( .A(v_length[24]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[24]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n180 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U232  ( .A(n5426), .B(n5672), .C(n5842), 
        .Y(\Decision_AXILiteS_s_axi_U/n655 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U231  ( .A(athresh[25]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[25]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n175 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U229  ( .A(v_length[25]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[25]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n177 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U228  ( .A(n5425), .B(n5671), .C(n5841), 
        .Y(\Decision_AXILiteS_s_axi_U/n654 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U227  ( .A(athresh[26]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[26]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n172 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U225  ( .A(v_length[26]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[26]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n174 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U224  ( .A(n5424), .B(n5670), .C(n5840), 
        .Y(\Decision_AXILiteS_s_axi_U/n653 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U223  ( .A(athresh[27]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[27]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n169 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U221  ( .A(v_length[27]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[27]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n171 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U220  ( .A(n5423), .B(n5669), .C(n5839), 
        .Y(\Decision_AXILiteS_s_axi_U/n652 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U219  ( .A(athresh[28]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[28]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n166 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U217  ( .A(v_length[28]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[28]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n168 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U216  ( .A(n5422), .B(n5668), .C(n5838), 
        .Y(\Decision_AXILiteS_s_axi_U/n651 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U215  ( .A(athresh[29]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[29]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n163 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U213  ( .A(v_length[29]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[29]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n165 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U212  ( .A(n5421), .B(n5667), .C(n5837), 
        .Y(\Decision_AXILiteS_s_axi_U/n650 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U211  ( .A(athresh[30]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[30]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n160 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U209  ( .A(v_length[30]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[30]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n162 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U208  ( .A(n5420), .B(n5666), .C(n5836), 
        .Y(\Decision_AXILiteS_s_axi_U/n649 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U207  ( .A(athresh[31]), .B(
        \Decision_AXILiteS_s_axi_U/n158 ), .C(vthresh[31]), .D(
        \Decision_AXILiteS_s_axi_U/n159 ), .Y(\Decision_AXILiteS_s_axi_U/n152 ) );
  AOI22X1 \Decision_AXILiteS_s_axi_U/U205  ( .A(v_length[31]), .B(
        \Decision_AXILiteS_s_axi_U/n155 ), .C(s_axi_AXILiteS_RDATA[31]), .D(
        n8918), .Y(\Decision_AXILiteS_s_axi_U/n154 ) );
  NAND3X1 \Decision_AXILiteS_s_axi_U/U204  ( .A(n5419), .B(n5665), .C(n5835), 
        .Y(\Decision_AXILiteS_s_axi_U/n648 ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[0]  ( .D(n4769), .CLK(n9115), 
        .Q(s_axi_AXILiteS_RDATA[0]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n692 ), .CLK(n9115), .Q(data[0]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[1]  ( .D(n4768), .CLK(n9115), 
        .Q(s_axi_AXILiteS_RDATA[1]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n691 ), .CLK(n9115), .Q(data[1]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[2]  ( .D(n4767), .CLK(n9115), 
        .Q(s_axi_AXILiteS_RDATA[2]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[2]  ( .D(
        \Decision_AXILiteS_s_axi_U/n690 ), .CLK(n9114), .Q(data[2]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[3]  ( .D(n4766), .CLK(n9114), 
        .Q(s_axi_AXILiteS_RDATA[3]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[3]  ( .D(
        \Decision_AXILiteS_s_axi_U/n689 ), .CLK(n9114), .Q(data[3]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[4]  ( .D(n9308), .CLK(n9114), 
        .Q(s_axi_AXILiteS_RDATA[4]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[4]  ( .D(
        \Decision_AXILiteS_s_axi_U/n688 ), .CLK(n9114), .Q(data[4]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[5]  ( .D(n9307), .CLK(n9114), 
        .Q(s_axi_AXILiteS_RDATA[5]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[5]  ( .D(
        \Decision_AXILiteS_s_axi_U/n687 ), .CLK(n9114), .Q(data[5]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[6]  ( .D(n9306), .CLK(n9114), 
        .Q(s_axi_AXILiteS_RDATA[6]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[6]  ( .D(
        \Decision_AXILiteS_s_axi_U/n686 ), .CLK(n9114), .Q(data[6]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[7]  ( .D(n4765), .CLK(n9114), 
        .Q(s_axi_AXILiteS_RDATA[7]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[7]  ( .D(
        \Decision_AXILiteS_s_axi_U/n685 ), .CLK(n9114), .Q(data[7]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[8]  ( .D(n4757), .CLK(n9114), 
        .Q(s_axi_AXILiteS_RDATA[8]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[8]  ( .D(
        \Decision_AXILiteS_s_axi_U/n684 ), .CLK(n9114), .Q(data[8]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[9]  ( .D(n4756), .CLK(n9113), 
        .Q(s_axi_AXILiteS_RDATA[9]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[9]  ( .D(
        \Decision_AXILiteS_s_axi_U/n683 ), .CLK(n9113), .Q(data[9]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[10]  ( .D(n4755), .CLK(n9113), 
        .Q(s_axi_AXILiteS_RDATA[10]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[10]  ( .D(
        \Decision_AXILiteS_s_axi_U/n682 ), .CLK(n9113), .Q(data[10]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[11]  ( .D(n4754), .CLK(n9113), 
        .Q(s_axi_AXILiteS_RDATA[11]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[11]  ( .D(
        \Decision_AXILiteS_s_axi_U/n681 ), .CLK(n9113), .Q(data[11]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[12]  ( .D(n4753), .CLK(n9113), 
        .Q(s_axi_AXILiteS_RDATA[12]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[12]  ( .D(
        \Decision_AXILiteS_s_axi_U/n680 ), .CLK(n9113), .Q(data[12]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[13]  ( .D(n4752), .CLK(n9113), 
        .Q(s_axi_AXILiteS_RDATA[13]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[13]  ( .D(
        \Decision_AXILiteS_s_axi_U/n679 ), .CLK(n9113), .Q(data[13]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[14]  ( .D(n4751), .CLK(n9113), 
        .Q(s_axi_AXILiteS_RDATA[14]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[14]  ( .D(
        \Decision_AXILiteS_s_axi_U/n678 ), .CLK(n9113), .Q(data[14]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[15]  ( .D(n4750), .CLK(n9113), 
        .Q(s_axi_AXILiteS_RDATA[15]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_data_reg[15]  ( .D(
        \Decision_AXILiteS_s_axi_U/n677 ), .CLK(n9112), .Q(data[15]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n724 ), .CLK(n9112), .Q(v_length[0]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n723 ), .CLK(n9112), .Q(v_length[1]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[2]  ( .D(
        \Decision_AXILiteS_s_axi_U/n722 ), .CLK(n9112), .Q(v_length[2]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[3]  ( .D(
        \Decision_AXILiteS_s_axi_U/n721 ), .CLK(n9112), .Q(v_length[3]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[4]  ( .D(
        \Decision_AXILiteS_s_axi_U/n720 ), .CLK(n9112), .Q(v_length[4]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[5]  ( .D(
        \Decision_AXILiteS_s_axi_U/n719 ), .CLK(n9112), .Q(v_length[5]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[6]  ( .D(
        \Decision_AXILiteS_s_axi_U/n718 ), .CLK(n9112), .Q(v_length[6]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[7]  ( .D(
        \Decision_AXILiteS_s_axi_U/n717 ), .CLK(n9112), .Q(v_length[7]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[8]  ( .D(
        \Decision_AXILiteS_s_axi_U/n716 ), .CLK(n9112), .Q(v_length[8]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[9]  ( .D(
        \Decision_AXILiteS_s_axi_U/n715 ), .CLK(n9112), .Q(v_length[9]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[10]  ( .D(
        \Decision_AXILiteS_s_axi_U/n714 ), .CLK(n9112), .Q(v_length[10]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[11]  ( .D(
        \Decision_AXILiteS_s_axi_U/n713 ), .CLK(n9112), .Q(v_length[11]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[12]  ( .D(
        \Decision_AXILiteS_s_axi_U/n712 ), .CLK(n9111), .Q(v_length[12]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[13]  ( .D(
        \Decision_AXILiteS_s_axi_U/n711 ), .CLK(n9111), .Q(v_length[13]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[14]  ( .D(
        \Decision_AXILiteS_s_axi_U/n710 ), .CLK(n9111), .Q(v_length[14]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[15]  ( .D(
        \Decision_AXILiteS_s_axi_U/n709 ), .CLK(n9111), .Q(v_length[15]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[16]  ( .D(n4749), .CLK(n9111), 
        .Q(s_axi_AXILiteS_RDATA[16]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[16]  ( .D(
        \Decision_AXILiteS_s_axi_U/n708 ), .CLK(n9111), .Q(v_length[16]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[17]  ( .D(n4748), .CLK(n9111), 
        .Q(s_axi_AXILiteS_RDATA[17]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[17]  ( .D(
        \Decision_AXILiteS_s_axi_U/n707 ), .CLK(n9111), .Q(v_length[17]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[18]  ( .D(n4747), .CLK(n9111), 
        .Q(s_axi_AXILiteS_RDATA[18]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[18]  ( .D(
        \Decision_AXILiteS_s_axi_U/n706 ), .CLK(n9111), .Q(v_length[18]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[19]  ( .D(n4746), .CLK(n9111), 
        .Q(s_axi_AXILiteS_RDATA[19]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[19]  ( .D(
        \Decision_AXILiteS_s_axi_U/n705 ), .CLK(n9111), .Q(v_length[19]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[20]  ( .D(n4745), .CLK(n9111), 
        .Q(s_axi_AXILiteS_RDATA[20]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[20]  ( .D(
        \Decision_AXILiteS_s_axi_U/n704 ), .CLK(n9110), .Q(v_length[20]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[21]  ( .D(n4744), .CLK(n9110), 
        .Q(s_axi_AXILiteS_RDATA[21]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[21]  ( .D(
        \Decision_AXILiteS_s_axi_U/n703 ), .CLK(n9110), .Q(v_length[21]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[22]  ( .D(n4743), .CLK(n9110), 
        .Q(s_axi_AXILiteS_RDATA[22]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[22]  ( .D(
        \Decision_AXILiteS_s_axi_U/n702 ), .CLK(n9110), .Q(v_length[22]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[23]  ( .D(n4742), .CLK(n9110), 
        .Q(s_axi_AXILiteS_RDATA[23]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[23]  ( .D(
        \Decision_AXILiteS_s_axi_U/n701 ), .CLK(n9110), .Q(v_length[23]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[24]  ( .D(n4741), .CLK(n9110), 
        .Q(s_axi_AXILiteS_RDATA[24]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[24]  ( .D(
        \Decision_AXILiteS_s_axi_U/n700 ), .CLK(n9110), .Q(v_length[24]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[25]  ( .D(n4740), .CLK(n9110), 
        .Q(s_axi_AXILiteS_RDATA[25]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[25]  ( .D(
        \Decision_AXILiteS_s_axi_U/n699 ), .CLK(n9110), .Q(v_length[25]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[26]  ( .D(n4739), .CLK(n9110), 
        .Q(s_axi_AXILiteS_RDATA[26]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[26]  ( .D(
        \Decision_AXILiteS_s_axi_U/n698 ), .CLK(n9110), .Q(v_length[26]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[27]  ( .D(n4738), .CLK(n9109), 
        .Q(s_axi_AXILiteS_RDATA[27]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[27]  ( .D(
        \Decision_AXILiteS_s_axi_U/n697 ), .CLK(n9109), .Q(v_length[27]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[28]  ( .D(n4737), .CLK(n9109), 
        .Q(s_axi_AXILiteS_RDATA[28]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[28]  ( .D(
        \Decision_AXILiteS_s_axi_U/n696 ), .CLK(n9109), .Q(v_length[28]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[29]  ( .D(n4736), .CLK(n9109), 
        .Q(s_axi_AXILiteS_RDATA[29]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[29]  ( .D(
        \Decision_AXILiteS_s_axi_U/n695 ), .CLK(n9109), .Q(v_length[29]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[30]  ( .D(n4735), .CLK(n9109), 
        .Q(s_axi_AXILiteS_RDATA[30]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[30]  ( .D(
        \Decision_AXILiteS_s_axi_U/n694 ), .CLK(n9109), .Q(v_length[30]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rdata_reg[31]  ( .D(n4734), .CLK(n9109), 
        .Q(s_axi_AXILiteS_RDATA[31]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_length_reg[31]  ( .D(
        \Decision_AXILiteS_s_axi_U/n693 ), .CLK(n9109), .Q(v_length[31]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n756 ), .CLK(n9109), .Q(a_length[0]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n755 ), .CLK(n9109), .Q(a_length[1]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[2]  ( .D(
        \Decision_AXILiteS_s_axi_U/n754 ), .CLK(n9109), .Q(a_length[2]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[3]  ( .D(
        \Decision_AXILiteS_s_axi_U/n753 ), .CLK(n9108), .Q(a_length[3]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[4]  ( .D(
        \Decision_AXILiteS_s_axi_U/n752 ), .CLK(n9108), .Q(a_length[4]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[5]  ( .D(
        \Decision_AXILiteS_s_axi_U/n751 ), .CLK(n9108), .Q(a_length[5]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[6]  ( .D(
        \Decision_AXILiteS_s_axi_U/n750 ), .CLK(n9108), .Q(a_length[6]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[7]  ( .D(
        \Decision_AXILiteS_s_axi_U/n749 ), .CLK(n9108), .Q(a_length[7]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[8]  ( .D(
        \Decision_AXILiteS_s_axi_U/n748 ), .CLK(n9108), .Q(a_length[8]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[9]  ( .D(
        \Decision_AXILiteS_s_axi_U/n747 ), .CLK(n9108), .Q(a_length[9]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[10]  ( .D(
        \Decision_AXILiteS_s_axi_U/n746 ), .CLK(n9108), .Q(a_length[10]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[11]  ( .D(
        \Decision_AXILiteS_s_axi_U/n745 ), .CLK(n9108), .Q(a_length[11]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[12]  ( .D(
        \Decision_AXILiteS_s_axi_U/n744 ), .CLK(n9108), .Q(a_length[12]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[13]  ( .D(
        \Decision_AXILiteS_s_axi_U/n743 ), .CLK(n9108), .Q(a_length[13]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[14]  ( .D(
        \Decision_AXILiteS_s_axi_U/n742 ), .CLK(n9108), .Q(a_length[14]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[15]  ( .D(
        \Decision_AXILiteS_s_axi_U/n741 ), .CLK(n9108), .Q(a_length[15]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[16]  ( .D(
        \Decision_AXILiteS_s_axi_U/n740 ), .CLK(n9107), .Q(a_length[16]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[17]  ( .D(
        \Decision_AXILiteS_s_axi_U/n739 ), .CLK(n9107), .Q(a_length[17]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[18]  ( .D(
        \Decision_AXILiteS_s_axi_U/n738 ), .CLK(n9107), .Q(a_length[18]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[19]  ( .D(
        \Decision_AXILiteS_s_axi_U/n737 ), .CLK(n9107), .Q(a_length[19]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[20]  ( .D(
        \Decision_AXILiteS_s_axi_U/n736 ), .CLK(n9107), .Q(a_length[20]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[21]  ( .D(
        \Decision_AXILiteS_s_axi_U/n735 ), .CLK(n9107), .Q(a_length[21]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[22]  ( .D(
        \Decision_AXILiteS_s_axi_U/n734 ), .CLK(n9107), .Q(a_length[22]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[23]  ( .D(
        \Decision_AXILiteS_s_axi_U/n733 ), .CLK(n9107), .Q(a_length[23]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[24]  ( .D(
        \Decision_AXILiteS_s_axi_U/n732 ), .CLK(n9107), .Q(a_length[24]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[25]  ( .D(
        \Decision_AXILiteS_s_axi_U/n731 ), .CLK(n9107), .Q(a_length[25]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[26]  ( .D(
        \Decision_AXILiteS_s_axi_U/n730 ), .CLK(n9107), .Q(a_length[26]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[27]  ( .D(
        \Decision_AXILiteS_s_axi_U/n729 ), .CLK(n9107), .Q(a_length[27]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[28]  ( .D(
        \Decision_AXILiteS_s_axi_U/n728 ), .CLK(n9107), .Q(a_length[28]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[29]  ( .D(
        \Decision_AXILiteS_s_axi_U/n727 ), .CLK(n9106), .Q(a_length[29]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[30]  ( .D(
        \Decision_AXILiteS_s_axi_U/n726 ), .CLK(n9106), .Q(a_length[30]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_length_reg[31]  ( .D(
        \Decision_AXILiteS_s_axi_U/n725 ), .CLK(n9106), .Q(a_length[31]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_flip_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n764 ), .CLK(n9106), .Q(v_flip[0]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_flip_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n763 ), .CLK(n9106), .Q(v_flip[1]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_flip_reg[2]  ( .D(
        \Decision_AXILiteS_s_axi_U/n762 ), .CLK(n9106), .Q(v_flip[2]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_flip_reg[3]  ( .D(
        \Decision_AXILiteS_s_axi_U/n761 ), .CLK(n9106), .Q(v_flip[3]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_flip_reg[4]  ( .D(
        \Decision_AXILiteS_s_axi_U/n760 ), .CLK(n9106), .Q(v_flip[4]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_flip_reg[5]  ( .D(
        \Decision_AXILiteS_s_axi_U/n759 ), .CLK(n9106), .Q(v_flip[5]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_flip_reg[6]  ( .D(
        \Decision_AXILiteS_s_axi_U/n758 ), .CLK(n9106), .Q(v_flip[6]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_v_flip_reg[7]  ( .D(
        \Decision_AXILiteS_s_axi_U/n757 ), .CLK(n9106), .Q(v_flip[7]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_flip_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n772 ), .CLK(n9106), .Q(a_flip[0]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_flip_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n771 ), .CLK(n9106), .Q(a_flip[1]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_flip_reg[2]  ( .D(
        \Decision_AXILiteS_s_axi_U/n770 ), .CLK(n9105), .Q(a_flip[2]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_flip_reg[3]  ( .D(
        \Decision_AXILiteS_s_axi_U/n769 ), .CLK(n9105), .Q(a_flip[3]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_flip_reg[4]  ( .D(
        \Decision_AXILiteS_s_axi_U/n768 ), .CLK(n9105), .Q(a_flip[4]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_flip_reg[5]  ( .D(
        \Decision_AXILiteS_s_axi_U/n767 ), .CLK(n9105), .Q(a_flip[5]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_flip_reg[6]  ( .D(
        \Decision_AXILiteS_s_axi_U/n766 ), .CLK(n9105), .Q(a_flip[6]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_a_flip_reg[7]  ( .D(
        \Decision_AXILiteS_s_axi_U/n765 ), .CLK(n9105), .Q(a_flip[7]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n804 ), .CLK(n9105), .Q(vthresh[0]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n803 ), .CLK(n9105), .Q(vthresh[1]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[2]  ( .D(
        \Decision_AXILiteS_s_axi_U/n802 ), .CLK(n9105), .Q(vthresh[2]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[3]  ( .D(
        \Decision_AXILiteS_s_axi_U/n801 ), .CLK(n9105), .Q(vthresh[3]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[4]  ( .D(
        \Decision_AXILiteS_s_axi_U/n800 ), .CLK(n9105), .Q(vthresh[4]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[5]  ( .D(
        \Decision_AXILiteS_s_axi_U/n799 ), .CLK(n9105), .Q(vthresh[5]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[6]  ( .D(
        \Decision_AXILiteS_s_axi_U/n798 ), .CLK(n9105), .Q(vthresh[6]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[7]  ( .D(
        \Decision_AXILiteS_s_axi_U/n797 ), .CLK(n9104), .Q(vthresh[7]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[8]  ( .D(
        \Decision_AXILiteS_s_axi_U/n796 ), .CLK(n9104), .Q(vthresh[8]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[9]  ( .D(
        \Decision_AXILiteS_s_axi_U/n795 ), .CLK(n9104), .Q(vthresh[9]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[10]  ( .D(
        \Decision_AXILiteS_s_axi_U/n794 ), .CLK(n9104), .Q(vthresh[10]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[11]  ( .D(
        \Decision_AXILiteS_s_axi_U/n793 ), .CLK(n9104), .Q(vthresh[11]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[12]  ( .D(
        \Decision_AXILiteS_s_axi_U/n792 ), .CLK(n9104), .Q(vthresh[12]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[13]  ( .D(
        \Decision_AXILiteS_s_axi_U/n791 ), .CLK(n9104), .Q(vthresh[13]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[14]  ( .D(
        \Decision_AXILiteS_s_axi_U/n790 ), .CLK(n9104), .Q(vthresh[14]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[15]  ( .D(
        \Decision_AXILiteS_s_axi_U/n789 ), .CLK(n9104), .Q(vthresh[15]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[16]  ( .D(
        \Decision_AXILiteS_s_axi_U/n788 ), .CLK(n9104), .Q(vthresh[16]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[17]  ( .D(
        \Decision_AXILiteS_s_axi_U/n787 ), .CLK(n9104), .Q(vthresh[17]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[18]  ( .D(
        \Decision_AXILiteS_s_axi_U/n786 ), .CLK(n9104), .Q(vthresh[18]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[19]  ( .D(
        \Decision_AXILiteS_s_axi_U/n785 ), .CLK(n9104), .Q(vthresh[19]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[20]  ( .D(
        \Decision_AXILiteS_s_axi_U/n784 ), .CLK(n9103), .Q(vthresh[20]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[21]  ( .D(
        \Decision_AXILiteS_s_axi_U/n783 ), .CLK(n9103), .Q(vthresh[21]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[22]  ( .D(
        \Decision_AXILiteS_s_axi_U/n782 ), .CLK(n9103), .Q(vthresh[22]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[23]  ( .D(
        \Decision_AXILiteS_s_axi_U/n781 ), .CLK(n9103), .Q(vthresh[23]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[24]  ( .D(
        \Decision_AXILiteS_s_axi_U/n780 ), .CLK(n9103), .Q(vthresh[24]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[25]  ( .D(
        \Decision_AXILiteS_s_axi_U/n779 ), .CLK(n9103), .Q(vthresh[25]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[26]  ( .D(
        \Decision_AXILiteS_s_axi_U/n778 ), .CLK(n9103), .Q(vthresh[26]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[27]  ( .D(
        \Decision_AXILiteS_s_axi_U/n777 ), .CLK(n9103), .Q(vthresh[27]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[28]  ( .D(
        \Decision_AXILiteS_s_axi_U/n776 ), .CLK(n9103), .Q(vthresh[28]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[29]  ( .D(
        \Decision_AXILiteS_s_axi_U/n775 ), .CLK(n9103), .Q(vthresh[29]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[30]  ( .D(
        \Decision_AXILiteS_s_axi_U/n774 ), .CLK(n9103), .Q(vthresh[30]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_vthresh_reg[31]  ( .D(
        \Decision_AXILiteS_s_axi_U/n773 ), .CLK(n9103), .Q(vthresh[31]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n836 ), .CLK(n9103), .Q(athresh[0]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n835 ), .CLK(n9102), .Q(athresh[1]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[2]  ( .D(
        \Decision_AXILiteS_s_axi_U/n834 ), .CLK(n9102), .Q(athresh[2]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[3]  ( .D(
        \Decision_AXILiteS_s_axi_U/n833 ), .CLK(n9102), .Q(athresh[3]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[4]  ( .D(
        \Decision_AXILiteS_s_axi_U/n832 ), .CLK(n9102), .Q(athresh[4]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[5]  ( .D(
        \Decision_AXILiteS_s_axi_U/n831 ), .CLK(n9102), .Q(athresh[5]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[6]  ( .D(
        \Decision_AXILiteS_s_axi_U/n830 ), .CLK(n9102), .Q(athresh[6]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[7]  ( .D(
        \Decision_AXILiteS_s_axi_U/n829 ), .CLK(n9102), .Q(athresh[7]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[8]  ( .D(
        \Decision_AXILiteS_s_axi_U/n828 ), .CLK(n9102), .Q(athresh[8]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[9]  ( .D(
        \Decision_AXILiteS_s_axi_U/n827 ), .CLK(n9102), .Q(athresh[9]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[10]  ( .D(
        \Decision_AXILiteS_s_axi_U/n826 ), .CLK(n9102), .Q(athresh[10]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[11]  ( .D(
        \Decision_AXILiteS_s_axi_U/n825 ), .CLK(n9102), .Q(athresh[11]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[12]  ( .D(
        \Decision_AXILiteS_s_axi_U/n824 ), .CLK(n9102), .Q(athresh[12]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[13]  ( .D(
        \Decision_AXILiteS_s_axi_U/n823 ), .CLK(n9102), .Q(athresh[13]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[14]  ( .D(
        \Decision_AXILiteS_s_axi_U/n822 ), .CLK(n9101), .Q(athresh[14]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[15]  ( .D(
        \Decision_AXILiteS_s_axi_U/n821 ), .CLK(n9101), .Q(athresh[15]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[16]  ( .D(
        \Decision_AXILiteS_s_axi_U/n820 ), .CLK(n9101), .Q(athresh[16]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[17]  ( .D(
        \Decision_AXILiteS_s_axi_U/n819 ), .CLK(n9101), .Q(athresh[17]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[18]  ( .D(
        \Decision_AXILiteS_s_axi_U/n818 ), .CLK(n9101), .Q(athresh[18]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[19]  ( .D(
        \Decision_AXILiteS_s_axi_U/n817 ), .CLK(n9101), .Q(athresh[19]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[20]  ( .D(
        \Decision_AXILiteS_s_axi_U/n816 ), .CLK(n9101), .Q(athresh[20]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[21]  ( .D(
        \Decision_AXILiteS_s_axi_U/n815 ), .CLK(n9101), .Q(athresh[21]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[22]  ( .D(
        \Decision_AXILiteS_s_axi_U/n814 ), .CLK(n9101), .Q(athresh[22]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[23]  ( .D(
        \Decision_AXILiteS_s_axi_U/n813 ), .CLK(n9101), .Q(athresh[23]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[24]  ( .D(
        \Decision_AXILiteS_s_axi_U/n812 ), .CLK(n9101), .Q(athresh[24]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[25]  ( .D(
        \Decision_AXILiteS_s_axi_U/n811 ), .CLK(n9101), .Q(athresh[25]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[26]  ( .D(
        \Decision_AXILiteS_s_axi_U/n810 ), .CLK(n9101), .Q(athresh[26]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[27]  ( .D(
        \Decision_AXILiteS_s_axi_U/n809 ), .CLK(n9100), .Q(athresh[27]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[28]  ( .D(
        \Decision_AXILiteS_s_axi_U/n808 ), .CLK(n9100), .Q(athresh[28]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[29]  ( .D(
        \Decision_AXILiteS_s_axi_U/n807 ), .CLK(n9100), .Q(athresh[29]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[30]  ( .D(
        \Decision_AXILiteS_s_axi_U/n806 ), .CLK(n9100), .Q(athresh[30]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_athresh_reg[31]  ( .D(
        \Decision_AXILiteS_s_axi_U/n805 ), .CLK(n9100), .Q(athresh[31]) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_reset_params_V_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n837 ), .CLK(n9100), .Q(\reset_params_V[0] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_reset_V_V_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n838 ), .CLK(n9100), .Q(\reset_V_V[0] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_reset_A_V_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n839 ), .CLK(n9100), .Q(\reset_A_V[0] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n840 ), .CLK(n9100), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[0] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n841 ), .CLK(n9100), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[1] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[2]  ( .D(
        \Decision_AXILiteS_s_axi_U/n842 ), .CLK(n9100), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[2] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[3]  ( .D(
        \Decision_AXILiteS_s_axi_U/n843 ), .CLK(n9100), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[3] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[4]  ( .D(
        \Decision_AXILiteS_s_axi_U/n844 ), .CLK(n9100), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[4] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[5]  ( .D(
        \Decision_AXILiteS_s_axi_U/n845 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[5] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[6]  ( .D(
        \Decision_AXILiteS_s_axi_U/n846 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[6] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[7]  ( .D(
        \Decision_AXILiteS_s_axi_U/n847 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[7] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[8]  ( .D(
        \Decision_AXILiteS_s_axi_U/n848 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[8] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[9]  ( .D(
        \Decision_AXILiteS_s_axi_U/n849 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[9] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[10]  ( .D(
        \Decision_AXILiteS_s_axi_U/n850 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[10] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[11]  ( .D(
        \Decision_AXILiteS_s_axi_U/n851 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[11] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[12]  ( .D(
        \Decision_AXILiteS_s_axi_U/n852 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[12] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[13]  ( .D(
        \Decision_AXILiteS_s_axi_U/n853 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[13] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[14]  ( .D(
        \Decision_AXILiteS_s_axi_U/n854 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[14] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_return_reg[15]  ( .D(
        \Decision_AXILiteS_s_axi_U/n855 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_ap_return[15] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_isr_reg[1]  ( .D(n4758), .CLK(n9099), 
        .Q(\Decision_AXILiteS_s_axi_U/int_isr[1] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_isr_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n857 ), .CLK(n9099), .Q(
        \Decision_AXILiteS_s_axi_U/int_isr[0] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ier_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n858 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/int_ier[0] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ier_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n859 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/int_ier[1] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_gie_reg  ( .D(
        \Decision_AXILiteS_s_axi_U/n860 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/int_gie ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_start_reg  ( .D(
        \Decision_AXILiteS_s_axi_U/n861 ), .CLK(n9098), .Q(ap_start) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_auto_restart_reg  ( .D(
        \Decision_AXILiteS_s_axi_U/n862 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/int_auto_restart ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/int_ap_done_reg  ( .D(n4770), .CLK(n9098), .Q(\Decision_AXILiteS_s_axi_U/int_ap_done ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/rstate_reg[0]  ( .D(n9275), .CLK(n9098), 
        .Q(\Decision_AXILiteS_s_axi_U/rstate[0] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/waddr_reg[0]  ( .D(
        \Decision_AXILiteS_s_axi_U/n865 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/waddr[0] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/waddr_reg[1]  ( .D(
        \Decision_AXILiteS_s_axi_U/n866 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/waddr[1] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/waddr_reg[2]  ( .D(
        \Decision_AXILiteS_s_axi_U/n867 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/waddr[2] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/waddr_reg[3]  ( .D(
        \Decision_AXILiteS_s_axi_U/n868 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/waddr[3] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/waddr_reg[4]  ( .D(
        \Decision_AXILiteS_s_axi_U/n869 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/waddr[4] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/waddr_reg[5]  ( .D(
        \Decision_AXILiteS_s_axi_U/n870 ), .CLK(n9098), .Q(
        \Decision_AXILiteS_s_axi_U/waddr[5] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/waddr_reg[6]  ( .D(
        \Decision_AXILiteS_s_axi_U/n871 ), .CLK(n9097), .Q(
        \Decision_AXILiteS_s_axi_U/waddr[6] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/wstate_reg[1]  ( .D(n9276), .CLK(n9097), 
        .Q(\Decision_AXILiteS_s_axi_U/wstate[1] ) );
  DFFPOSX1 \Decision_AXILiteS_s_axi_U/wstate_reg[0]  ( .D(n4762), .CLK(n9097), 
        .Q(\Decision_AXILiteS_s_axi_U/wstate[0] ) );
  NOR3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1221  ( 
        .A(n9822), .B(n9823), .C(n9809), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n14 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1217  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11045), .C(n8208), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1228 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1214  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11044), .C(n7966), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1227 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1211  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11043), .C(n7749), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1226 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1208  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11042), .C(n7551), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1225 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1205  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11041), .C(n7370), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1224 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1202  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11040), .C(n7207), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1223 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1199  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11039), .C(n7053), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1222 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1196  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11038), .C(n6912), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1221 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1193  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11037), .C(n6778), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1220 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1190  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11036), .C(n6657), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1219 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1187  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11035), .C(n7369), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1218 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1184  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11034), .C(n7206), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1217 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1181  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11033), .C(n7052), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1216 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1178  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11032), .C(n6911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1215 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1175  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11031), .C(n6546), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1214 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1172  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), .B(n11030), .C(n6435), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1213 )
         );
  NOR3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1170  ( 
        .A(n9822), .B(n8888), .C(n9809), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n13 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1167  ( 
        .A(n9793), .B(n8917), .C(n8207), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1212 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1164  ( 
        .A(n9794), .B(n8917), .C(n7965), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1211 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1161  ( 
        .A(n9795), .B(n8917), .C(n7748), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1210 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1158  ( 
        .A(n9796), .B(n8917), .C(n7550), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1209 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1155  ( 
        .A(n9797), .B(n8917), .C(n7368), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1208 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1152  ( 
        .A(n9798), .B(n8917), .C(n7205), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1207 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1149  ( 
        .A(n9799), .B(n8917), .C(n7051), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1206 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1146  ( 
        .A(n9800), .B(n8917), .C(n6910), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1205 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1143  ( 
        .A(n9801), .B(n8917), .C(n6777), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1204 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1140  ( 
        .A(n9802), .B(n8917), .C(n6656), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1203 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1137  ( 
        .A(n9803), .B(n8917), .C(n6545), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1202 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1134  ( 
        .A(n9804), .B(n8917), .C(n6434), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1201 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1131  ( 
        .A(n9805), .B(n8917), .C(n6326), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1200 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1128  ( 
        .A(n9806), .B(n8917), .C(n6232), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1199 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1125  ( 
        .A(n9807), .B(n8917), .C(n7747), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1198 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1122  ( 
        .A(n9808), .B(n8917), .C(n7549), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1197 )
         );
  NOR3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1121  ( 
        .A(n9823), .B(n8889), .C(n9809), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n15 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1118  ( 
        .A(n9793), .B(n8916), .C(n7964), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1196 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1116  ( 
        .A(n9794), .B(n8916), .C(n8206), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1195 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1114  ( 
        .A(n9795), .B(n8916), .C(n7548), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1194 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1112  ( 
        .A(n9796), .B(n8916), .C(n7746), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1193 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1110  ( 
        .A(n9797), .B(n8916), .C(n7204), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1192 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1108  ( 
        .A(n9798), .B(n8916), .C(n7367), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1191 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1106  ( 
        .A(n9799), .B(n8916), .C(n6909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1190 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1104  ( 
        .A(n9800), .B(n8916), .C(n7050), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1189 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1102  ( 
        .A(n9801), .B(n8916), .C(n6655), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1188 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1100  ( 
        .A(n9802), .B(n8916), .C(n6776), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1187 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1098  ( 
        .A(n9803), .B(n8916), .C(n6433), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1186 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1096  ( 
        .A(n9804), .B(n8916), .C(n6544), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1185 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1094  ( 
        .A(n9805), .B(n8916), .C(n6231), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1184 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1092  ( 
        .A(n9806), .B(n8916), .C(n6325), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1183 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1090  ( 
        .A(n9807), .B(n8916), .C(n7547), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1182 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1088  ( 
        .A(n9808), .B(n8916), .C(n7745), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1181 )
         );
  NOR3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1087  ( 
        .A(n8888), .B(n8889), .C(n9809), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n17 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1084  ( 
        .A(n9793), .B(n8915), .C(n7744), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1180 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1082  ( 
        .A(n9794), .B(n8915), .C(n7546), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1179 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1080  ( 
        .A(n9795), .B(n8915), .C(n8205), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1178 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1078  ( 
        .A(n9796), .B(n8915), .C(n7963), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1177 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1076  ( 
        .A(n9797), .B(n8915), .C(n7049), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1176 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1074  ( 
        .A(n9798), .B(n8915), .C(n6908), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1175 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1072  ( 
        .A(n9799), .B(n8915), .C(n7366), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1174 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1070  ( 
        .A(n9800), .B(n8915), .C(n7203), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1173 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1068  ( 
        .A(n9801), .B(n8915), .C(n6543), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1172 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1066  ( 
        .A(n9802), .B(n8915), .C(n6432), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1171 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1064  ( 
        .A(n9803), .B(n8915), .C(n6775), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1170 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1062  ( 
        .A(n9804), .B(n8915), .C(n6654), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1169 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1060  ( 
        .A(n9805), .B(n8915), .C(n6150), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1168 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1058  ( 
        .A(n9806), .B(n8915), .C(n6083), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1167 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1056  ( 
        .A(n9807), .B(n8915), .C(n8204), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1166 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1054  ( 
        .A(n9808), .B(n8915), .C(n7962), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1165 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1050  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 ), .C(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n688 ), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n807 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1046  ( 
        .A(n9466), .B(n11029), .C(n7961), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1164 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1043  ( 
        .A(n9466), .B(n11028), .C(n8203), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1163 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1040  ( 
        .A(n9466), .B(n11027), .C(n7545), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1162 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1037  ( 
        .A(n9466), .B(n11026), .C(n7743), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1161 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1034  ( 
        .A(n9466), .B(n11025), .C(n7202), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1160 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1031  ( 
        .A(n9466), .B(n11024), .C(n7365), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1159 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1028  ( 
        .A(n9466), .B(n11023), .C(n6907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1158 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1025  ( 
        .A(n9466), .B(n11022), .C(n7048), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1157 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1022  ( 
        .A(n9466), .B(n11021), .C(n6653), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1156 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1019  ( 
        .A(n9466), .B(n11020), .C(n6774), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1155 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1016  ( 
        .A(n9466), .B(n11019), .C(n7201), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1154 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1013  ( 
        .A(n9466), .B(n11018), .C(n7364), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1153 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1010  ( 
        .A(n9466), .B(n11017), .C(n6906), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1152 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1007  ( 
        .A(n9466), .B(n11016), .C(n7047), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1151 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1004  ( 
        .A(n9466), .B(n11015), .C(n6431), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1150 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U1001  ( 
        .A(n9466), .B(n11014), .C(n6542), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1149 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U998  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 ), .C(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n669 ), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n757 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U996  ( 
        .A(n9793), .B(n8913), .C(n7544), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1148 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U994  ( 
        .A(n9794), .B(n8913), .C(n7742), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1147 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U992  ( 
        .A(n9795), .B(n8913), .C(n7960), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1146 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U990  ( 
        .A(n9796), .B(n8913), .C(n8202), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1145 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U988  ( 
        .A(n9797), .B(n8913), .C(n6905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1144 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U986  ( 
        .A(n9798), .B(n8913), .C(n7046), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1143 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U984  ( 
        .A(n9799), .B(n8913), .C(n7200), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1142 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U982  ( 
        .A(n9800), .B(n8913), .C(n7363), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1141 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U980  ( 
        .A(n9801), .B(n8913), .C(n6430), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1140 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U978  ( 
        .A(n9802), .B(n8913), .C(n6541), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1139 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U976  ( 
        .A(n9803), .B(n8913), .C(n6652), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1138 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U974  ( 
        .A(n9804), .B(n8913), .C(n6773), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1137 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U972  ( 
        .A(n9805), .B(n8913), .C(n6082), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1136 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U970  ( 
        .A(n9806), .B(n8913), .C(n6149), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1135 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U968  ( 
        .A(n9807), .B(n8913), .C(n7959), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1134 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U966  ( 
        .A(n9808), .B(n8913), .C(n8201), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1133 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U964  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 ), .C(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n688 ), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n740 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U962  ( 
        .A(n9793), .B(n8911), .C(n7362), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1132 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U960  ( 
        .A(n9794), .B(n8911), .C(n7199), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1131 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U958  ( 
        .A(n9795), .B(n8911), .C(n7045), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1130 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U956  ( 
        .A(n9796), .B(n8911), .C(n6904), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1129 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U954  ( 
        .A(n9797), .B(n8911), .C(n8200), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1128 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U952  ( 
        .A(n9798), .B(n8911), .C(n7958), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1127 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U950  ( 
        .A(n9799), .B(n8911), .C(n7741), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1126 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U948  ( 
        .A(n9800), .B(n8911), .C(n7543), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1125 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U946  ( 
        .A(n9801), .B(n8911), .C(n6324), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1124 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U944  ( 
        .A(n9802), .B(n8911), .C(n6230), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1123 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U942  ( 
        .A(n9803), .B(n8911), .C(n6148), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1122 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U940  ( 
        .A(n9804), .B(n8911), .C(n6081), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1121 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U938  ( 
        .A(n9805), .B(n8911), .C(n6772), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1120 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U936  ( 
        .A(n9806), .B(n8911), .C(n6651), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1119 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U934  ( 
        .A(n9807), .B(n8911), .C(n7044), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1118 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U932  ( 
        .A(n9808), .B(n8911), .C(n6903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1117 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U931  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 ), .C(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n669 ), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n723 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U929  ( 
        .A(n9793), .B(n8909), .C(n7198), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1116 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U927  ( 
        .A(n9794), .B(n8909), .C(n7361), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1115 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U925  ( 
        .A(n9795), .B(n8909), .C(n6902), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1114 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U923  ( 
        .A(n9796), .B(n8909), .C(n7043), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1113 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U921  ( 
        .A(n9797), .B(n8909), .C(n7957), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1112 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U919  ( 
        .A(n9798), .B(n8909), .C(n8199), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1111 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U917  ( 
        .A(n9799), .B(n8909), .C(n7542), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1110 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U915  ( 
        .A(n9800), .B(n8909), .C(n7740), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1109 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U913  ( 
        .A(n9801), .B(n8909), .C(n6229), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1108 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U911  ( 
        .A(n9802), .B(n8909), .C(n6323), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1107 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U909  ( 
        .A(n9803), .B(n8909), .C(n6080), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1106 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U907  ( 
        .A(n9804), .B(n8909), .C(n6147), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1105 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U905  ( 
        .A(n9805), .B(n8909), .C(n6650), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1104 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U903  ( 
        .A(n9806), .B(n8909), .C(n6771), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1103 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U901  ( 
        .A(n9807), .B(n8909), .C(n6901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1102 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U899  ( 
        .A(n9808), .B(n8909), .C(n7042), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1101 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U898  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n670 ), .B(n8889), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n688 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n706 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U896  ( 
        .A(n9793), .B(n8907), .C(n7041), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1100 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U894  ( 
        .A(n9794), .B(n8907), .C(n6900), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1099 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U892  ( 
        .A(n9795), .B(n8907), .C(n7360), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1098 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U890  ( 
        .A(n9796), .B(n8907), .C(n7197), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1097 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U888  ( 
        .A(n9797), .B(n8907), .C(n7739), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1096 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U886  ( 
        .A(n9798), .B(n8907), .C(n7541), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1095 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U884  ( 
        .A(n9799), .B(n8907), .C(n8198), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1094 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U882  ( 
        .A(n9800), .B(n8907), .C(n7956), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1093 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U880  ( 
        .A(n9801), .B(n8907), .C(n6146), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1092 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U878  ( 
        .A(n9802), .B(n8907), .C(n6079), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1091 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U876  ( 
        .A(n9803), .B(n8907), .C(n6322), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1090 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U874  ( 
        .A(n9804), .B(n8907), .C(n6228), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1089 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U872  ( 
        .A(n9805), .B(n8907), .C(n6540), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1088 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U870  ( 
        .A(n9806), .B(n8907), .C(n6429), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1087 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U868  ( 
        .A(n9807), .B(n8907), .C(n7359), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1086 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U866  ( 
        .A(n9808), .B(n8907), .C(n7196), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1085 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U865  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n669 ), .B(n8889), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n670 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n689 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U863  ( 
        .A(n9793), .B(n8905), .C(n6899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1084 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U861  ( 
        .A(n9794), .B(n8905), .C(n7040), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1083 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U859  ( 
        .A(n9795), .B(n8905), .C(n7195), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1082 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U857  ( 
        .A(n9796), .B(n8905), .C(n7358), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1081 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U855  ( 
        .A(n9797), .B(n8905), .C(n7540), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1080 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U853  ( 
        .A(n9798), .B(n8905), .C(n7738), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1079 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U851  ( 
        .A(n9799), .B(n8905), .C(n7955), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1078 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U849  ( 
        .A(n9800), .B(n8905), .C(n8197), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1077 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U847  ( 
        .A(n9801), .B(n8905), .C(n6078), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1076 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U845  ( 
        .A(n9802), .B(n8905), .C(n6145), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1075 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U843  ( 
        .A(n9803), .B(n8905), .C(n6227), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1074 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U841  ( 
        .A(n9804), .B(n8905), .C(n6321), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1073 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U839  ( 
        .A(n9805), .B(n8905), .C(n6428), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1072 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U837  ( 
        .A(n9806), .B(n8905), .C(n6539), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1071 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U835  ( 
        .A(n9807), .B(n8905), .C(n7194), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1070 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U833  ( 
        .A(n9808), .B(n8905), .C(n7357), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1069 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U832  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n670 ), .B(n9822), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n688 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n671 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U830  ( 
        .A(n9793), .B(n8903), .C(n6770), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1068 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U828  ( 
        .A(n9794), .B(n8903), .C(n6649), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1067 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U826  ( 
        .A(n9795), .B(n8903), .C(n6538), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1066 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U824  ( 
        .A(n9796), .B(n8903), .C(n6427), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1065 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U822  ( 
        .A(n9797), .B(n8903), .C(n6320), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1064 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U820  ( 
        .A(n9798), .B(n8903), .C(n6226), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1063 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U818  ( 
        .A(n9799), .B(n8903), .C(n6144), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1062 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U816  ( 
        .A(n9800), .B(n8903), .C(n6077), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1061 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U814  ( 
        .A(n9801), .B(n8903), .C(n8196), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1060 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U812  ( 
        .A(n9802), .B(n8903), .C(n7954), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1059 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U810  ( 
        .A(n9803), .B(n8903), .C(n7737), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1058 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U808  ( 
        .A(n9804), .B(n8903), .C(n7539), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1057 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U806  ( 
        .A(n9805), .B(n8903), .C(n7356), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1056 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U804  ( 
        .A(n9806), .B(n8903), .C(n7193), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1055 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U802  ( 
        .A(n9807), .B(n8903), .C(n6537), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1054 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U800  ( 
        .A(n9808), .B(n8903), .C(n6426), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1053 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U799  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n669 ), .B(n9822), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n670 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n652 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U797  ( 
        .A(n9793), .B(n8901), .C(n6648), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1052 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U795  ( 
        .A(n9794), .B(n8901), .C(n6769), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1051 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U793  ( 
        .A(n9795), .B(n8901), .C(n6425), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1050 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U791  ( 
        .A(n9796), .B(n8901), .C(n6536), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1049 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U789  ( 
        .A(n9797), .B(n8901), .C(n6225), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1048 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U787  ( 
        .A(n9798), .B(n8901), .C(n6319), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1047 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U785  ( 
        .A(n9799), .B(n8901), .C(n6076), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1046 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U783  ( 
        .A(n9800), .B(n8901), .C(n6143), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1045 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U781  ( 
        .A(n9801), .B(n8901), .C(n7953), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1044 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U779  ( 
        .A(n9802), .B(n8901), .C(n8195), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1043 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U777  ( 
        .A(n9803), .B(n8901), .C(n7538), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1042 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U775  ( 
        .A(n9804), .B(n8901), .C(n7736), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1041 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U773  ( 
        .A(n9805), .B(n8901), .C(n7192), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1040 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U771  ( 
        .A(n9806), .B(n8901), .C(n7355), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1039 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U769  ( 
        .A(n9807), .B(n8901), .C(n6424), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1038 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U767  ( 
        .A(n9808), .B(n8901), .C(n6535), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1037 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U766  ( 
        .A(n4693), .B(n9809), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n650 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U764  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 ), .B(n8888), .C(n9470), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n649 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U760  ( 
        .A(n9469), .B(n11013), .C(n7735), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1036 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U757  ( 
        .A(n9469), .B(n11012), .C(n7537), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1035 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U754  ( 
        .A(n9469), .B(n11011), .C(n8194), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1034 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U751  ( 
        .A(n9469), .B(n11010), .C(n7952), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1033 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U748  ( 
        .A(n9469), .B(n11009), .C(n7039), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1032 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U745  ( 
        .A(n9469), .B(n11008), .C(n6898), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1031 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U742  ( 
        .A(n9469), .B(n11007), .C(n7354), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1030 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U739  ( 
        .A(n9469), .B(n11006), .C(n7191), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1029 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U736  ( 
        .A(n9469), .B(n11005), .C(n6534), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1028 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U733  ( 
        .A(n9469), .B(n11004), .C(n6423), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1027 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U730  ( 
        .A(n9469), .B(n11003), .C(n7038), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1026 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U727  ( 
        .A(n9469), .B(n11002), .C(n6897), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1025 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U724  ( 
        .A(n9469), .B(n11001), .C(n7353), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1024 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U721  ( 
        .A(n9469), .B(n11000), .C(n7190), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1023 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U718  ( 
        .A(n9469), .B(n10999), .C(n6768), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1022 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U715  ( 
        .A(n9469), .B(n10998), .C(n6647), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1021 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U714  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 ), .B(n9823), .C(n9470), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n615 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U710  ( 
        .A(n9468), .B(n10997), .C(n7536), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1020 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U707  ( 
        .A(n9468), .B(n10996), .C(n7734), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1019 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U704  ( 
        .A(n9468), .B(n10995), .C(n7951), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1018 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U701  ( 
        .A(n9468), .B(n10994), .C(n8193), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1017 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U698  ( 
        .A(n9468), .B(n10993), .C(n6896), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1016 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U695  ( 
        .A(n9468), .B(n10992), .C(n7037), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1015 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U692  ( 
        .A(n9468), .B(n10991), .C(n7189), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1014 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U689  ( 
        .A(n9468), .B(n10990), .C(n7352), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1013 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U686  ( 
        .A(n9468), .B(n10989), .C(n6422), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1012 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U683  ( 
        .A(n9468), .B(n10988), .C(n6533), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1011 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U680  ( 
        .A(n9468), .B(n10987), .C(n6895), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1010 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U677  ( 
        .A(n9468), .B(n10986), .C(n7036), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1009 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U674  ( 
        .A(n9468), .B(n10985), .C(n7188), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1008 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U671  ( 
        .A(n9468), .B(n10984), .C(n7351), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1007 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U668  ( 
        .A(n9468), .B(n10983), .C(n6646), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1006 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U665  ( 
        .A(n9468), .B(n10982), .C(n6767), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1005 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U664  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 ), .B(n8888), .C(n9470), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n550 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U662  ( 
        .A(n9793), .B(n8899), .C(n6532), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1004 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U660  ( 
        .A(n9794), .B(n8899), .C(n6421), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1003 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U658  ( 
        .A(n9795), .B(n8899), .C(n6766), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1002 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U656  ( 
        .A(n9796), .B(n8899), .C(n6645), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1001 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U654  ( 
        .A(n9797), .B(n8899), .C(n6142), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1000 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U652  ( 
        .A(n9798), .B(n8899), .C(n6075), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n999 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U650  ( 
        .A(n9799), .B(n8899), .C(n6318), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n998 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U648  ( 
        .A(n9800), .B(n8899), .C(n6224), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n997 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U646  ( 
        .A(n9801), .B(n8899), .C(n7733), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n996 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U644  ( 
        .A(n9802), .B(n8899), .C(n7535), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n995 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U642  ( 
        .A(n9803), .B(n8899), .C(n8192), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n994 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U640  ( 
        .A(n9804), .B(n8899), .C(n7950), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n993 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U638  ( 
        .A(n9805), .B(n8899), .C(n7035), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n992 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U636  ( 
        .A(n9806), .B(n8899), .C(n6894), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n991 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U634  ( 
        .A(n9807), .B(n8899), .C(n6765), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n990 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U632  ( 
        .A(n9808), .B(n8899), .C(n6644), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n989 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U631  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 ), .B(n9823), .C(n9470), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n547 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U627  ( 
        .A(n9467), .B(n10981), .C(n7350), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n988 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U624  ( 
        .A(n9467), .B(n10980), .C(n7187), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n987 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U621  ( 
        .A(n9467), .B(n10979), .C(n7034), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n986 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U618  ( 
        .A(n9467), .B(n10978), .C(n6893), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n985 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U615  ( 
        .A(n9467), .B(n10977), .C(n8191), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n984 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U612  ( 
        .A(n9467), .B(n10976), .C(n7949), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n983 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U609  ( 
        .A(n9467), .B(n10975), .C(n7732), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n982 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U606  ( 
        .A(n9467), .B(n10974), .C(n7534), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n981 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U603  ( 
        .A(n9467), .B(n10973), .C(n6317), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n980 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U600  ( 
        .A(n9467), .B(n10972), .C(n6223), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n979 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U597  ( 
        .A(n9467), .B(n10971), .C(n8190), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n978 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U594  ( 
        .A(n9467), .B(n10970), .C(n7948), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n977 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U591  ( 
        .A(n9467), .B(n10969), .C(n7731), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n976 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U588  ( 
        .A(n9467), .B(n10968), .C(n7533), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n975 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U585  ( 
        .A(n9467), .B(n10967), .C(n6141), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n974 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U582  ( 
        .A(n9467), .B(n10966), .C(n6074), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n973 )
         );
  NOR3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U581  ( 
        .A(n6019), .B(n5971), .C(n6012), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n411 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U580  ( 
        .A(n8889), .B(n8888), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n411 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n513 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U575  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10965), .C(n7186), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n972 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U572  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10964), .C(n7349), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n971 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U569  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10963), .C(n6892), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n970 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U566  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10962), .C(n7033), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n969 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U563  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10961), .C(n7947), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n968 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U560  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10960), .C(n8189), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n967 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U557  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10959), .C(n7532), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n966 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U554  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10958), .C(n7730), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n965 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U551  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10957), .C(n6222), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n964 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U548  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10956), .C(n6316), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n963 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U545  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10955), .C(n7946), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n962 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U542  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10954), .C(n8188), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n961 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U539  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10953), .C(n7531), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n960 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U536  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10952), .C(n7729), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n959 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U533  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10951), .C(n6073), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n958 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U530  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), .B(n10950), .C(n6140), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n957 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U529  ( 
        .A(n8889), .B(n9823), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n411 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n479 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U524  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10949), .C(n7032), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n956 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U521  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10948), .C(n6891), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n955 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U518  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10947), .C(n7348), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n954 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U515  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10946), .C(n7185), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n953 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U512  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10945), .C(n7728), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n952 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U509  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10944), .C(n7530), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n951 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U506  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10943), .C(n8187), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n950 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U503  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10942), .C(n7945), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n949 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U500  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10941), .C(n6139), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n948 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U497  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10940), .C(n6072), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n947 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U494  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10939), .C(n7727), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n946 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U491  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10938), .C(n7529), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n945 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U488  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10937), .C(n8186), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n944 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U485  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10936), .C(n7944), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n943 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U482  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10935), .C(n6315), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n942 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U479  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), .B(n10934), .C(n6221), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n941 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U478  ( 
        .A(n8888), .B(n9822), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n411 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n445 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U473  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10933), .C(n6890), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n940 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U470  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10932), .C(n7031), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n939 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U467  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10931), .C(n7184), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n938 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U464  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10930), .C(n7347), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n937 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U461  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10929), .C(n7528), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n936 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U458  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10928), .C(n7726), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n935 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U455  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10927), .C(n7943), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n934 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U452  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10926), .C(n8185), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n933 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U449  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10925), .C(n6071), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n932 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U446  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10924), .C(n6138), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n931 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U443  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10923), .C(n7527), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n930 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U440  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10922), .C(n7725), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n929 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U437  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10921), .C(n7942), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n928 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U434  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10920), .C(n8184), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n927 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U431  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10919), .C(n6220), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n926 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U428  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), .B(n10918), .C(n6314), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n925 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U427  ( 
        .A(n9823), .B(n9822), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n411 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n410 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U422  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10917), .C(n6764), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n924 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U419  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10916), .C(n6643), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n923 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U416  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10915), .C(n6531), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n922 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U413  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10914), .C(n6420), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n921 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U410  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10913), .C(n6313), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n920 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U407  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10912), .C(n6219), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n919 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U404  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10911), .C(n6137), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n918 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U401  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10910), .C(n6070), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n917 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U398  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10909), .C(n8183), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n916 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U395  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10908), .C(n7941), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n915 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U392  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10907), .C(n6312), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n914 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U389  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10906), .C(n6218), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n913 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U386  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10905), .C(n6136), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n912 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U383  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10904), .C(n6069), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n911 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U380  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10903), .C(n7724), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n910 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U377  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), .B(n10902), .C(n7526), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n909 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U374  ( 
        .A(n9823), .B(n9822), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n362 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n375 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U372  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n362 ), .B(n9822), .C(n8888), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n373 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U370  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][15] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][15] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n367 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U369  ( 
        .A(n9823), .B(n4693), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n372 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U366  ( 
        .A(n8888), .B(n4693), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n371 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U364  ( 
        .A(n9823), .B(n4693), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n370 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U362  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][15] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][15] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n369 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U361  ( 
        .A(n5418), .B(n5664), .C(n5834), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n355 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U360  ( 
        .A(n8888), .B(n4693), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n365 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U358  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n362 ), .B(n9823), .C(n8889), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n363 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U356  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][15] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][15] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n357 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U355  ( 
        .A(n8888), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n362 ), 
        .C(n8889), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n361 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U350  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][15] ), .B(n8866), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][15] ), .D(n8864), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n359 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U349  ( 
        .A(n5417), .B(n5663), .C(n5833), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n356 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U345  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][15] ), .B(n8862), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][15] ), .D(n8860), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n349 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U343  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][15] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][15] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n351 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U342  ( 
        .A(n5416), .B(n5662), .C(n5832), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n344 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U341  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][15] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][15] ), .D(n8876), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n346 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U339  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][15] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][15] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n348 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U338  ( 
        .A(n5415), .B(n5661), .C(n5831), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n345 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U334  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n342 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n343 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n340 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U332  ( 
        .A(n5499), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n340 ), 
        .C(n5892), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n908 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U330  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][14] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][14] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n336 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U328  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][14] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][14] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n338 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U327  ( 
        .A(n5414), .B(n5660), .C(n5830), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n331 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U326  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][14] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][14] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n333 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U324  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][14] ), .B(n8866), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][14] ), .D(n8864), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n335 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U323  ( 
        .A(n5413), .B(n5659), .C(n5829), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n332 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U321  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][14] ), .B(n8862), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][14] ), .D(n8860), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n328 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U319  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][14] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][14] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n330 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U318  ( 
        .A(n5412), .B(n5658), .C(n5828), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n323 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U317  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][14] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][14] ), .D(n8876), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n325 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U315  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][14] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][14] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n327 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U314  ( 
        .A(n5411), .B(n5657), .C(n5827), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n324 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U312  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n321 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n322 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n319 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U310  ( 
        .A(n5498), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n319 ), 
        .C(n5891), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n907 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U308  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][13] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][13] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n315 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U306  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][13] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][13] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n317 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U305  ( 
        .A(n5410), .B(n5656), .C(n5826), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n310 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U304  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][13] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][13] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n312 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U302  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][13] ), .B(n8866), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][13] ), .D(n8864), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n314 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U301  ( 
        .A(n5409), .B(n5655), .C(n5825), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n311 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U299  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][13] ), .B(n8862), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][13] ), .D(n8860), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n307 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U297  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][13] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][13] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n309 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U296  ( 
        .A(n5408), .B(n5654), .C(n5824), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n302 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U295  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][13] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][13] ), .D(n8876), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n304 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U293  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][13] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][13] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n306 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U292  ( 
        .A(n5407), .B(n5653), .C(n5823), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n303 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U290  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n300 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n301 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n298 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U288  ( 
        .A(n5497), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n298 ), 
        .C(n5890), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n906 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U286  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][12] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][12] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n294 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U284  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][12] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][12] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n296 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U283  ( 
        .A(n5406), .B(n5652), .C(n5822), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n289 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U282  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][12] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][12] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n291 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U280  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][12] ), .B(n8866), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][12] ), .D(n8864), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n293 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U279  ( 
        .A(n5405), .B(n5651), .C(n5821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n290 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U277  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][12] ), .B(n8862), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][12] ), .D(n8860), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n286 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U275  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][12] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][12] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n288 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U274  ( 
        .A(n5404), .B(n5650), .C(n5820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n281 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U273  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][12] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][12] ), .D(n8876), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n283 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U271  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][12] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][12] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n285 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U270  ( 
        .A(n5403), .B(n5649), .C(n5819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n282 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U268  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n279 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n280 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n277 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U266  ( 
        .A(n5496), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n277 ), 
        .C(n5889), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n905 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U264  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][11] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][11] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n273 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U262  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][11] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][11] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n275 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U261  ( 
        .A(n5402), .B(n5648), .C(n5818), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n268 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U260  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][11] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][11] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n270 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U258  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][11] ), .B(n8866), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][11] ), .D(n8864), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n272 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U257  ( 
        .A(n5401), .B(n5647), .C(n5817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n269 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U255  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][11] ), .B(n8862), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][11] ), .D(n8860), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n265 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U253  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][11] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][11] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n267 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U252  ( 
        .A(n5400), .B(n5646), .C(n5816), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n260 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U251  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][11] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][11] ), .D(n8876), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n262 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U249  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][11] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][11] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n264 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U248  ( 
        .A(n5399), .B(n5645), .C(n5815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n261 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U246  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n258 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n259 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n256 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U244  ( 
        .A(n5495), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n256 ), 
        .C(n5888), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n904 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U242  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][10] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][10] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n252 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U240  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][10] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][10] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n254 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U239  ( 
        .A(n5398), .B(n5644), .C(n5814), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n247 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U238  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][10] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][10] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n249 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U236  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][10] ), .B(n8866), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][10] ), .D(n8864), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n251 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U235  ( 
        .A(n5397), .B(n5643), .C(n5813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n248 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U233  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][10] ), .B(n8862), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][10] ), .D(n8860), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n244 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U231  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][10] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][10] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n246 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U230  ( 
        .A(n5396), .B(n5642), .C(n5812), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n239 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U229  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][10] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][10] ), .D(n8876), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n241 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U227  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][10] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][10] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n243 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U226  ( 
        .A(n5395), .B(n5641), .C(n5811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n240 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U224  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n237 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n238 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n235 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U222  ( 
        .A(n5494), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n235 ), 
        .C(n5887), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n903 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U220  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][9] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][9] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n231 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U218  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][9] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][9] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n233 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U217  ( 
        .A(n5394), .B(n5640), .C(n5810), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n226 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U216  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][9] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][9] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n228 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U214  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][9] ), .B(n8866), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][9] ), .D(n8864), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n230 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U213  ( 
        .A(n5393), .B(n5639), .C(n5809), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n227 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U211  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][9] ), .B(n8862), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][9] ), .D(n8860), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n223 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U209  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][9] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][9] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n225 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U208  ( 
        .A(n5392), .B(n5638), .C(n5808), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n218 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U207  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][9] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][9] ), .D(n8876), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n220 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U205  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][9] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][9] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n222 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U204  ( 
        .A(n5391), .B(n5637), .C(n5807), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n219 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U202  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n216 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n217 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n214 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U200  ( 
        .A(n5493), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n214 ), 
        .C(n5886), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n902 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U198  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][8] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][8] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n210 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U196  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][8] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][8] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n212 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U195  ( 
        .A(n5390), .B(n5636), .C(n5806), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n205 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U194  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][8] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][8] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n207 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U192  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][8] ), .B(n8866), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][8] ), .D(n8864), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n209 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U191  ( 
        .A(n5389), .B(n5635), .C(n5805), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n206 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U189  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][8] ), .B(n8862), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][8] ), .D(n8860), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n202 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U187  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][8] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][8] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n204 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U186  ( 
        .A(n5388), .B(n5634), .C(n5804), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n197 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U185  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][8] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][8] ), .D(n8876), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n199 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U183  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][8] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][8] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n201 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U182  ( 
        .A(n5387), .B(n5633), .C(n5803), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n198 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U180  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n195 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n196 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n193 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U178  ( 
        .A(n5492), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n193 ), 
        .C(n5885), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n901 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U176  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][7] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][7] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n189 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U174  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][7] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][7] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n191 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U173  ( 
        .A(n5386), .B(n5632), .C(n5802), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n184 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U172  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][7] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][7] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n186 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U170  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][7] ), .B(n8867), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][7] ), .D(n8865), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n188 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U169  ( 
        .A(n5385), .B(n5631), .C(n5801), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n185 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U167  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][7] ), .B(n8863), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][7] ), .D(n8861), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n181 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U165  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][7] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][7] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n183 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U164  ( 
        .A(n5384), .B(n5630), .C(n5800), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n176 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U163  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][7] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][7] ), .D(n8877), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n178 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U161  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][7] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][7] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n180 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U160  ( 
        .A(n5383), .B(n5629), .C(n5799), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n177 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U158  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n174 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n175 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n172 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U156  ( 
        .A(n5491), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n172 ), 
        .C(n5884), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n900 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U154  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][6] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][6] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n168 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U152  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][6] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][6] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n170 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U151  ( 
        .A(n5382), .B(n5628), .C(n5798), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n163 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U150  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][6] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][6] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n165 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U148  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][6] ), .B(n8867), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][6] ), .D(n8865), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n167 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U147  ( 
        .A(n5381), .B(n5627), .C(n5797), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n164 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U145  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][6] ), .B(n8863), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][6] ), .D(n8861), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n160 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U143  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][6] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][6] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n162 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U142  ( 
        .A(n5380), .B(n5626), .C(n5796), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n155 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U141  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][6] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][6] ), .D(n8877), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n157 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U139  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][6] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][6] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n159 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U138  ( 
        .A(n5379), .B(n5625), .C(n5795), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n156 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U136  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n153 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n154 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n151 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U134  ( 
        .A(n5490), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n151 ), 
        .C(n5883), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n899 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U132  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][5] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][5] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n147 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U130  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][5] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][5] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n149 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U129  ( 
        .A(n5378), .B(n5624), .C(n5794), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n142 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U128  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][5] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][5] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n144 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U126  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][5] ), .B(n8867), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][5] ), .D(n8865), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n146 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U125  ( 
        .A(n5377), .B(n5623), .C(n5793), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n143 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U123  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][5] ), .B(n8863), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][5] ), .D(n8861), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n139 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U121  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][5] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][5] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n141 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U120  ( 
        .A(n5376), .B(n5622), .C(n5792), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n134 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U119  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][5] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][5] ), .D(n8877), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n136 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U117  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][5] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][5] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n138 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U116  ( 
        .A(n5375), .B(n5621), .C(n5791), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n135 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U114  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n132 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n133 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n130 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U112  ( 
        .A(n5489), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n130 ), 
        .C(n5882), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n898 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U110  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][4] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][4] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n126 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U108  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][4] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][4] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n128 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U107  ( 
        .A(n5374), .B(n5620), .C(n5790), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n121 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U106  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][4] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][4] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n123 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U104  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][4] ), .B(n8867), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][4] ), .D(n8865), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n125 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U103  ( 
        .A(n5373), .B(n5619), .C(n5789), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n122 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U101  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][4] ), .B(n8863), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][4] ), .D(n8861), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n118 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U99  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][4] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][4] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n120 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U98  ( 
        .A(n5372), .B(n5618), .C(n5788), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n113 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U97  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][4] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][4] ), .D(n8877), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n115 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U95  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][4] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][4] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n117 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U94  ( 
        .A(n5371), .B(n5617), .C(n5787), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n114 )
         );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U92  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n111 ), .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n112 ), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n109 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U90  ( 
        .A(n5488), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n109 ), 
        .C(n5881), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n897 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U88  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][3] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][3] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n105 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U86  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][3] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][3] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n107 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U85  ( 
        .A(n5370), .B(n5616), .C(n5786), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n100 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U84  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][3] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][3] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n102 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U82  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][3] ), .B(n8867), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][3] ), .D(n8865), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n104 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U81  ( 
        .A(n5369), .B(n5615), .C(n5785), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n101 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U79  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][3] ), .B(n8863), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][3] ), .D(n8861), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n97 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U77  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][3] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][3] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n99 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U76  ( 
        .A(n5368), .B(n5614), .C(n5784), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n92 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U75  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][3] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][3] ), .D(n8877), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n94 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U73  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][3] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][3] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n96 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U72  ( 
        .A(n5367), .B(n5613), .C(n5783), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n93 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U70  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n90 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n91 ), 
        .C(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n88 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U68  ( 
        .A(n5487), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n88 ), 
        .C(n5880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n896 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U66  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][2] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][2] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n84 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U64  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][2] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][2] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n86 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U63  ( 
        .A(n5366), .B(n5612), .C(n5782), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n79 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U62  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][2] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][2] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n81 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U60  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][2] ), .B(n8867), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][2] ), .D(n8865), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n83 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U59  ( 
        .A(n5365), .B(n5611), .C(n5781), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n80 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U57  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][2] ), .B(n8863), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][2] ), .D(n8861), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n76 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U55  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][2] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][2] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n78 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U54  ( 
        .A(n5364), .B(n5610), .C(n5780), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n71 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U53  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][2] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][2] ), .D(n8877), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n73 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U51  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][2] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][2] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n75 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U50  ( 
        .A(n5363), .B(n5609), .C(n5779), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n72 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U48  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n69 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n70 ), 
        .C(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n67 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U46  ( 
        .A(n5486), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n67 ), 
        .C(n5879), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n895 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U44  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][1] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][1] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n63 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U42  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][1] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][1] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n65 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U41  ( 
        .A(n5362), .B(n5608), .C(n5778), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n58 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U40  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][1] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][1] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n60 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U38  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][1] ), .B(n8867), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][1] ), .D(n8865), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n62 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U37  ( 
        .A(n5361), .B(n5607), .C(n5777), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n59 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U35  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][1] ), .B(n8863), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][1] ), .D(n8861), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n55 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U33  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][1] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][1] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n57 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U32  ( 
        .A(n5360), .B(n5606), .C(n5776), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n50 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U31  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][1] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][1] ), .D(n8877), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n52 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U29  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][1] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][1] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n54 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U28  ( 
        .A(n5359), .B(n5605), .C(n5775), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n51 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U26  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n48 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n49 ), 
        .C(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n46 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U24  ( 
        .A(n5485), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n46 ), 
        .C(n5878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n894 )
         );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U22  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][0] ), .B(n9818), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][0] ), .D(n9819), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n36 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U20  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][0] ), .B(n9816), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][0] ), .D(n9815), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n38 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U19  ( 
        .A(n5358), .B(n5604), .C(n5774), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n26 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U18  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][0] ), .B(n9814), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][0] ), .D(n9820), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n28 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U16  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][0] ), .B(n8867), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][0] ), .D(n8865), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n30 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U15  ( 
        .A(n5357), .B(n5603), .C(n5773), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n27 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U13  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][0] ), .B(n8863), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][0] ), .D(n8861), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n18 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U11  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][0] ), .B(n9812), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][0] ), .D(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n20 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U10  ( 
        .A(n5356), .B(n5602), .C(n5772), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n8 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U9  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][0] ), .B(n9810), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][0] ), .D(n8877), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n10 ) );
  AOI22X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U7  ( 
        .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][0] ), .B(n8879), .C(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][0] ), .D(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n12 ) );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U6  ( 
        .A(n5355), .B(n5601), .C(n5771), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n9 ) );
  OAI21X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U4  ( 
        .A(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n5 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n6 ), 
        .C(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n2 )
         );
  NAND3X1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/U2  ( 
        .A(n5484), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n2 ), 
        .C(n5877), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n893 )
         );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[0]  ( 
        .D(n4718), .CLK(n9097), .Q(recentdatapoints_data_q0[0]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[1]  ( 
        .D(n4719), .CLK(n9097), .Q(recentdatapoints_data_q0[1]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[2]  ( 
        .D(n4720), .CLK(n9097), .Q(recentdatapoints_data_q0[2]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[3]  ( 
        .D(n4721), .CLK(n9097), .Q(recentdatapoints_data_q0[3]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[4]  ( 
        .D(n4722), .CLK(n9097), .Q(recentdatapoints_data_q0[4]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[5]  ( 
        .D(n4723), .CLK(n9097), .Q(recentdatapoints_data_q0[5]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[6]  ( 
        .D(n4724), .CLK(n9097), .Q(recentdatapoints_data_q0[6]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[7]  ( 
        .D(n4725), .CLK(n9097), .Q(recentdatapoints_data_q0[7]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[8]  ( 
        .D(n4726), .CLK(n9097), .Q(recentdatapoints_data_q0[8]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[9]  ( 
        .D(n4727), .CLK(n9097), .Q(recentdatapoints_data_q0[9]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[10]  ( 
        .D(n4728), .CLK(n9096), .Q(recentdatapoints_data_q0[10]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[11]  ( 
        .D(n4729), .CLK(n9096), .Q(recentdatapoints_data_q0[11]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[12]  ( 
        .D(n4730), .CLK(n9096), .Q(recentdatapoints_data_q0[12]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[13]  ( 
        .D(n4731), .CLK(n9096), .Q(recentdatapoints_data_q0[13]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[14]  ( 
        .D(n4732), .CLK(n9096), .Q(recentdatapoints_data_q0[14]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/q0_reg[15]  ( 
        .D(n4733), .CLK(n9096), .Q(recentdatapoints_data_q0[15]) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][0]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n909 ), .CLK(n9096), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][1]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n910 ), .CLK(n9096), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][2]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n911 ), .CLK(n9096), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][3]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n912 ), .CLK(n9096), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][4]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n913 ), .CLK(n9096), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][5]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n914 ), .CLK(n9096), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][6]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n915 ), .CLK(n9096), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][7]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n916 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][8]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n917 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][9]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n918 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][10]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n919 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][11]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n920 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][12]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n921 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][13]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n922 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][14]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n923 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[0][15]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n924 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][0]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n925 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][1]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n926 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][2]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n927 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][3]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n928 ), .CLK(n9095), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][4]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n929 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][5]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n930 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][6]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n931 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][7]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n932 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][8]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n933 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][9]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n934 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][10]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n935 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][11]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n936 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][12]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n937 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][13]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n938 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][14]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n939 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[1][15]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n940 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][0]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n941 ), .CLK(n9094), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][1]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n942 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][2]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n943 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][3]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n944 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][4]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n945 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][5]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n946 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][6]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n947 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][7]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n948 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][8]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n949 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][9]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n950 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][10]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n951 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][11]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n952 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][12]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n953 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][13]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n954 ), .CLK(n9093), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][14]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n955 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[2][15]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n956 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][0]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n957 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][1]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n958 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][2]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n959 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][3]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n960 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][4]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n961 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][5]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n962 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][6]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n963 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][7]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n964 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][8]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n965 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][9]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n966 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][10]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n967 ), .CLK(n9092), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][11]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n968 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][12]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n969 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][13]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n970 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][14]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n971 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[3][15]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n972 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][0]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n973 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][1]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n974 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][2]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n975 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][3]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n976 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][4]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n977 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][5]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n978 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][6]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n979 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][7]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n980 ), .CLK(n9091), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][8]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n981 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][9]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n982 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][10]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n983 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][11]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n984 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][12]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n985 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][13]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n986 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][14]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n987 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[4][15]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n988 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][0]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n989 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][1]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n990 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][2]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n991 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][3]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n992 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][4]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n993 ), .CLK(n9090), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][5]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n994 ), .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][6]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n995 ), .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][7]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n996 ), .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][8]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n997 ), .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][9]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n998 ), .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][10]  ( 
        .D(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n999 ), .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1000 ), 
        .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1001 ), 
        .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1002 ), 
        .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1003 ), 
        .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[5][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1004 ), 
        .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1005 ), 
        .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1006 ), 
        .CLK(n9089), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1007 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1008 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1009 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1010 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1011 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1012 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1013 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1014 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1015 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1016 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1017 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1018 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1019 ), 
        .CLK(n9088), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[6][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1020 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1021 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1022 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1023 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1024 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1025 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1026 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1027 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1028 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1029 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1030 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1031 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1032 ), 
        .CLK(n9087), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1033 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1034 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1035 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[7][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1036 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1037 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1038 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1039 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1040 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1041 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1042 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1043 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1044 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1045 ), 
        .CLK(n9086), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1046 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1047 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1048 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1049 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1050 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1051 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[8][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1052 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1053 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1054 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1055 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1056 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1057 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1058 ), 
        .CLK(n9085), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1059 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1060 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1061 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1062 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1063 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1064 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1065 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1066 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1067 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[9][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1068 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1069 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1070 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1071 ), 
        .CLK(n9084), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1072 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1073 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1074 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1075 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1076 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1077 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1078 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1079 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1080 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1081 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1082 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1083 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[10][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1084 ), 
        .CLK(n9083), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1085 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1086 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1087 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1088 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1089 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1090 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1091 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1092 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1093 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1094 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1095 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1096 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1097 ), 
        .CLK(n9082), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1098 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1099 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[11][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1100 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1101 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1102 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1103 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1104 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1105 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1106 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1107 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1108 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1109 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1110 ), 
        .CLK(n9081), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1111 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1112 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1113 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1114 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1115 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[12][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1116 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1117 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1118 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1119 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1120 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1121 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1122 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1123 ), 
        .CLK(n9080), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1124 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1125 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1126 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1127 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1128 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1129 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1130 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1131 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[13][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1132 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1133 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1134 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1135 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1136 ), 
        .CLK(n9079), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1137 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1138 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1139 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1140 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1141 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1142 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1143 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1144 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1145 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1146 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1147 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[14][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1148 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1149 ), 
        .CLK(n9078), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1150 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1151 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1152 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1153 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1154 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1155 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1156 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1157 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1158 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1159 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1160 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1161 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1162 ), 
        .CLK(n9077), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1163 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[15][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1164 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1165 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1166 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1167 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1168 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1169 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1170 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1171 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1172 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1173 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1174 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1175 ), 
        .CLK(n9076), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1176 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1177 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1178 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1179 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[16][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1180 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1181 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1182 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1183 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1184 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1185 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1186 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1187 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1188 ), 
        .CLK(n9075), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1189 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1190 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1191 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1192 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1193 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1194 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1195 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[17][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1196 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1197 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1198 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1199 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1200 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1201 ), 
        .CLK(n9074), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1202 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1203 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1204 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1205 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1206 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1207 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1208 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1209 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1210 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1211 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[18][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1212 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][15] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][0]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1213 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][0] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][1]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1214 ), 
        .CLK(n9073), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][1] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][2]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1215 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][2] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][3]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1216 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][3] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][4]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1217 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][4] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][5]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1218 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][5] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][6]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1219 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][6] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][7]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1220 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][7] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][8]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1221 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][8] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][9]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1222 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][9] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][10]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1223 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][10] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][11]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1224 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][11] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][12]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1225 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][12] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][13]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1226 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][13] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][14]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1227 ), 
        .CLK(n9072), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][14] ) );
  DFFPOSX1 \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram_reg[19][15]  ( 
        .D(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1228 ), 
        .CLK(n9071), .Q(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][15] ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U165  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ), .S(
        n9996), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n161 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U164  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ), .S(
        n9996), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n162 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U163  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ), .S(
        n9996), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n158 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U162  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ), .S(
        n9996), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n159 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U161  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ), .S(
        n9996), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n155 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U160  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n156 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U159  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n152 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U158  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n153 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U157  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n149 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U156  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n150 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U155  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n146 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U154  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n147 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U153  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n142 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U152  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n143 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U151  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n161 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n162 ), .S(n9995), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n160 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U150  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n158 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n159 ), .S(n9995), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n157 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U149  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n155 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n156 ), .S(n9995), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n154 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U148  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n152 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n153 ), .S(n9995), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n151 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U147  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n149 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n150 ), .S(n9995), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n148 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U146  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n146 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n147 ), .S(n9995), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n145 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U144  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n142 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n143 ), .S(n9995), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n141 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U143  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ), 
        .S(n9996), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n140 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U142  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ), .S(
        n8886), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n138 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U141  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ), .S(
        n8886), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n139 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U140  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ), .S(
        n8886), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n135 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U139  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ), .S(
        n8886), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n136 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U138  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ), .S(
        n8886), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n132 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U137  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ), 
        .S(n8886), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n133 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U136  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ), 
        .S(n8886), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n129 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U135  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ), 
        .S(n8886), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n130 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U134  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ), 
        .S(n8886), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n126 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U133  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ), 
        .S(n8887), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n127 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U132  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ), 
        .S(n8887), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n123 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U131  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ), 
        .S(n8887), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n124 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U130  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ), 
        .S(n8887), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n119 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U129  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ), 
        .S(n8887), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n120 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U128  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n138 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n139 ), .S(
        recentVBools_data_address0[1]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n137 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U127  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n135 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n136 ), .S(
        recentVBools_data_address0[1]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n134 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U126  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n132 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n133 ), .S(
        recentVBools_data_address0[1]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n131 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U125  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n129 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n130 ), .S(
        recentVBools_data_address0[1]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n128 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U124  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n126 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n127 ), .S(
        recentVBools_data_address0[1]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n125 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U123  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n123 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n124 ), .S(
        recentVBools_data_address0[1]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n122 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U121  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n119 ), .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n120 ), .S(
        recentVBools_data_address0[1]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n118 ) );
  MUX2X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U120  ( .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ), 
        .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ), 
        .S(n8887), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n117 ) );
  NAND3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U118  ( .A(
        n8413), .B(n8644), .C(n8887), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n44 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U113  ( .A(
        n8118), .B(n6027), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n83 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U112  ( .A(
        n8118), .B(n7101), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n83 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n116 ) );
  NAND3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U110  ( .A(
        recentVBools_data_address0[0]), .B(n8644), .C(n8413), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n42 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U109  ( .A(
        n7868), .B(n6027), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n82 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U108  ( .A(
        n7868), .B(n7101), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n82 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n115 ) );
  NAND3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U106  ( .A(
        n8887), .B(recentVBools_data_address0[2]), .C(
        recentVBools_data_address0[1]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n40 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U105  ( .A(
        n7867), .B(n6027), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n81 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U104  ( .A(
        n7867), .B(n7101), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n81 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n114 ) );
  NAND3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U103  ( .A(
        recentVBools_data_address0[0]), .B(recentVBools_data_address0[2]), .C(
        recentVBools_data_address0[1]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n38 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U102  ( .A(
        n8117), .B(n6027), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n80 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U101  ( .A(
        n8117), .B(n7101), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n80 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n113 ) );
  NAND3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U100  ( .A(
        n8644), .B(recentVBools_data_address0[2]), .C(n8887), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n36 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U99  ( .A(
        n7654), .B(n6027), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n79 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U98  ( .A(
        n7654), .B(n7101), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n79 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n112 ) );
  NAND3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U97  ( .A(
        n8644), .B(recentVBools_data_address0[2]), .C(
        recentVBools_data_address0[0]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n32 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U96  ( .A(
        n7270), .B(n6027), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n76 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U95  ( .A(
        n7270), .B(n7101), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n76 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n111 ) );
  NAND3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U91  ( .A(
        n6017), .B(recentVBools_data_address0[3]), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n18 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n64 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U88  ( .A(
        n7266), .B(n8875), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n73 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U87  ( .A(
        n7266), .B(n6035), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n73 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n110 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U85  ( .A(
        n7647), .B(n8875), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n70 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U84  ( .A(
        n7647), .B(n6035), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n70 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n109 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U83  ( .A(
        n8118), .B(n8875), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n69 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U82  ( .A(
        n8118), .B(n6035), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n69 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n108 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U81  ( .A(
        n7868), .B(n8875), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n68 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U80  ( .A(
        n7868), .B(n6035), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n68 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n107 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U79  ( .A(
        n7867), .B(n8875), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n67 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U78  ( .A(
        n7867), .B(n6035), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n67 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n106 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U77  ( .A(
        n8117), .B(n8875), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n66 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U76  ( .A(
        n8117), .B(n6035), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n66 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n105 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U75  ( .A(
        n7654), .B(n8875), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n65 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U74  ( .A(
        n7654), .B(n6035), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n65 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n104 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U73  ( .A(
        n7270), .B(n8875), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n63 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U72  ( .A(
        n7270), .B(n6035), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n63 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n103 ) );
  NAND3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U70  ( .A(
        n8108), .B(recentVBools_data_address0[4]), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n18 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n53 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U67  ( .A(
        n7266), .B(n8874), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n60 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U66  ( .A(
        n7266), .B(n6034), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n60 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n102 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U65  ( .A(
        n7647), .B(n8874), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n59 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U64  ( .A(
        n7647), .B(n6034), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n59 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n101 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U63  ( .A(
        n8118), .B(n8874), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n58 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U62  ( .A(
        n8118), .B(n6034), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n58 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n100 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U61  ( .A(
        n7868), .B(n8874), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n57 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U60  ( .A(
        n7868), .B(n6034), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n57 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n99 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U59  ( .A(
        n7867), .B(n8874), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n56 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U58  ( .A(
        n7867), .B(n6034), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n56 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n98 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U57  ( .A(
        n8117), .B(n8874), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n55 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U56  ( .A(
        n8117), .B(n6034), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n55 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n97 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U55  ( .A(
        n7654), .B(n8874), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n54 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U54  ( .A(
        n7654), .B(n6034), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n54 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n96 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U53  ( .A(
        n7270), .B(n8874), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n52 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U52  ( .A(
        n7270), .B(n6034), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n52 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n95 ) );
  NAND3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U51  ( .A(
        recentVBools_data_address0[3]), .B(recentVBools_data_address0[4]), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n18 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n35 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U48  ( .A(
        n8873), .B(n7266), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n49 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U47  ( .A(
        n7449), .B(n7266), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n49 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n94 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U46  ( .A(
        n8873), .B(n7647), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n47 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U45  ( .A(
        n7449), .B(n7647), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n47 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n93 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U44  ( .A(
        n8873), .B(n8118), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n45 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U43  ( .A(
        n7449), .B(n8118), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n45 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n92 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U42  ( .A(
        n8873), .B(n7868), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n43 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U41  ( .A(
        n7449), .B(n7868), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n43 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n91 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U40  ( .A(
        n8873), .B(n7867), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n41 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U39  ( .A(
        n7449), .B(n7867), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n41 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n90 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U38  ( .A(
        n8873), .B(n8117), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n39 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U37  ( .A(
        n7449), .B(n8117), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n39 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n89 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U36  ( .A(
        n8873), .B(n7654), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n37 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U35  ( .A(
        n7449), .B(n7654), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n37 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n88 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U34  ( .A(
        n8873), .B(n7270), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n34 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U33  ( .A(
        n7270), .B(n7449), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n34 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n87 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U31  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n137 ), .B(
        recentVBools_data_address0[2]), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n134 ), .D(n8413), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n29 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U30  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n131 ), .B(
        recentVBools_data_address0[2]), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n128 ), .D(n8413), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n31 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U28  ( .A(
        n8108), .B(n6934), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n30 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n21 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U27  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n125 ), .B(
        recentVBools_data_address0[2]), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n122 ), .D(n8413), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n24 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U26  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n118 ), .B(
        recentVBools_data_address0[2]), .C(n7405), .D(n8413), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n26 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U24  ( .A(
        n8108), .B(n7081), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n25 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n23 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U23  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n21 ), .B(
        recentVBools_data_address0[4]), .C(n6017), .D(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n23 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n20 ) );
  NOR3X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U22  ( .A(N466), 
        .B(n8981), .C(n5903), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n19 ) );
  AOI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U21  ( .A(
        \tmp_s_reg_1578[0] ), .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n18 ), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n19 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n15 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U17  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n160 ), .B(n8396), .C(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n157 ), .D(n9994), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n12 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U16  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n154 ), .B(n8396), .C(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n151 ), .D(n9994), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n14 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U13  ( .A(
        n9993), .B(n5698), .C(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n13 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n4 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U11  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n148 ), .B(n8396), .C(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n145 ), .D(n9994), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n7 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U10  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n141 ), .B(n8396), .C(n7795), .D(n9994), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n9 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U8  ( .A(n9993), .B(n5697), .C(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n8 ), 
        .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n6 ) );
  AOI22X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U7  ( .A(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n4 ), .B(n7630), 
        .C(n9992), .D(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n6 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n1 ) );
  OAI21X1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/U4  ( .A(n5530), .B(n10056), .C(n4938), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n85 ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/q1_reg[0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n85 ), .CLK(
        n9071), .Q(\recentVBools_data_q1[0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/q0_reg[0]  ( 
        .D(n4764), .CLK(n9071), .Q(\recentVBools_data_q0[0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[0][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n87 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[1][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n88 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[2][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n89 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[3][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n90 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[4][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n91 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[5][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n92 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[6][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n93 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[7][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n94 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[8][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n95 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[9][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n96 ), .CLK(
        n9071), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[10][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n97 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[11][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n98 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[12][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n99 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[13][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n100 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[14][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n101 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[15][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n102 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[16][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n103 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[17][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n104 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[18][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n105 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[19][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n106 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[20][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n107 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[21][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n108 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[22][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n109 ), .CLK(
        n9070), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[23][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n110 ), .CLK(
        n9069), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[24][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n111 ), .CLK(
        n9069), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[25][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n112 ), .CLK(
        n9069), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[26][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n113 ), .CLK(
        n9069), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[27][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n114 ), .CLK(
        n9069), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[28][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n115 ), .CLK(
        n9069), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ) );
  DFFPOSX1 \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram_reg[29][0]  ( 
        .D(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n116 ), .CLK(
        n9069), .Q(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U165  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ), .S(
        n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n160 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U164  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ), .S(
        n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n161 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U163  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ), .S(
        n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n157 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U162  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ), .S(
        n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n158 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U161  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ), .S(
        n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n154 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U160  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n155 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U159  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n151 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U158  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n152 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U157  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n148 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U156  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n149 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U155  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n145 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U154  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n146 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U153  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n142 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U152  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n143 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U151  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ), 
        .S(n10278), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n162 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U150  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n160 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n161 ), .S(
        n10277), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n159 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U149  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n157 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n158 ), .S(
        n10277), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n156 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U148  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n154 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n155 ), .S(
        n10277), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n153 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U147  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n151 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n152 ), .S(
        n10277), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n150 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U146  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n148 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n149 ), .S(
        n10277), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n147 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U145  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n145 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n146 ), .S(
        n10277), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n144 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U144  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n142 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n143 ), .S(
        n10277), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n141 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U143  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ), .S(
        n8884), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n138 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U142  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ), .S(
        n8884), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n139 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U141  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ), .S(
        n8884), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n135 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U140  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ), .S(
        n8884), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n136 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U139  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ), .S(
        n8884), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n132 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U138  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ), 
        .S(n8884), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n133 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U137  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ), 
        .S(n8884), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n129 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U136  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ), 
        .S(n8884), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n130 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U135  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ), 
        .S(n8884), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n126 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U134  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ), 
        .S(n8885), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n127 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U133  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ), 
        .S(n8885), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n123 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U132  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ), 
        .S(n8885), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n124 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U131  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ), 
        .S(n8885), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n120 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U130  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ), 
        .S(n8885), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n121 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U129  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ), 
        .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ), 
        .S(n8885), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n140 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U128  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n138 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n139 ), .S(
        recentABools_data_address0[1]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n137 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U127  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n135 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n136 ), .S(
        recentABools_data_address0[1]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n134 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U126  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n132 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n133 ), .S(
        recentABools_data_address0[1]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n131 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U125  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n129 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n130 ), .S(
        recentABools_data_address0[1]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n128 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U124  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n126 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n127 ), .S(
        recentABools_data_address0[1]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n125 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U123  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n123 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n124 ), .S(
        recentABools_data_address0[1]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n122 ) );
  MUX2X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U122  ( .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n120 ), .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n121 ), .S(
        recentABools_data_address0[1]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n119 ) );
  NAND3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U120  ( .A(
        n7648), .B(n8645), .C(n8885), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n46 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U115  ( .A(
        n6031), .B(n6024), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n85 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U114  ( .A(
        n6031), .B(n7267), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n85 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n118 ) );
  NAND3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U112  ( .A(
        recentABools_data_address0[0]), .B(n8645), .C(n7648), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n44 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U111  ( .A(
        n6030), .B(n6024), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n84 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U110  ( .A(
        n6030), .B(n7267), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n84 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n117 ) );
  NAND3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U108  ( .A(
        n8885), .B(recentABools_data_address0[2]), .C(
        recentABools_data_address0[1]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n42 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U107  ( .A(
        n8416), .B(n6024), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n83 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U106  ( .A(
        n8416), .B(n7267), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n83 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n116 ) );
  NAND3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U105  ( .A(
        recentABools_data_address0[0]), .B(recentABools_data_address0[2]), .C(
        recentABools_data_address0[1]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n40 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U104  ( .A(
        n8119), .B(n6024), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n82 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U103  ( .A(
        n8119), .B(n7267), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n82 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n115 ) );
  NAND3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U102  ( .A(
        n8645), .B(recentABools_data_address0[2]), .C(n8885), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n38 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U101  ( .A(
        n7869), .B(n6024), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n81 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U100  ( .A(
        n7869), .B(n7267), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n81 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n114 ) );
  NAND3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U99  ( .A(
        n8645), .B(recentABools_data_address0[2]), .C(
        recentABools_data_address0[0]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n34 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U98  ( .A(
        n7448), .B(n6024), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n78 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U97  ( .A(
        n7448), .B(n7267), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n78 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n113 ) );
  NAND3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U93  ( .A(
        n6016), .B(recentABools_data_address0[3]), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n19 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n66 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U90  ( .A(
        n7444), .B(n8872), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n75 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U89  ( .A(
        n7444), .B(n6033), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n75 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n112 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U87  ( .A(
        n6023), .B(n8872), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n72 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U86  ( .A(
        n6023), .B(n6033), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n72 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n111 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U85  ( .A(
        n6031), .B(n8872), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n71 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U84  ( .A(
        n6031), .B(n6033), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n71 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n110 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U83  ( .A(
        n6030), .B(n8872), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n70 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U82  ( .A(
        n6030), .B(n6033), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n70 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n109 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U81  ( .A(
        n8416), .B(n8872), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n69 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U80  ( .A(
        n8416), .B(n6033), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n69 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n108 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U79  ( .A(
        n8119), .B(n8872), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n68 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U78  ( .A(
        n8119), .B(n6033), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n68 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n107 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U77  ( .A(
        n7869), .B(n8872), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n67 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U76  ( .A(
        n7869), .B(n6033), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n67 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n106 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U75  ( .A(
        n7448), .B(n8872), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n65 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U74  ( .A(
        n7448), .B(n6033), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n65 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n105 ) );
  NAND3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U72  ( .A(
        n8402), .B(recentABools_data_address0[4]), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n19 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n55 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U69  ( .A(
        n7444), .B(n8871), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n62 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U68  ( .A(
        n7444), .B(n6032), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n62 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n104 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U67  ( .A(
        n6023), .B(n8871), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n61 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U66  ( .A(
        n6023), .B(n6032), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n61 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n103 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U65  ( .A(
        n6031), .B(n8871), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n60 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U64  ( .A(
        n6031), .B(n6032), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n60 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n102 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U63  ( .A(
        n6030), .B(n8871), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n59 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U62  ( .A(
        n6030), .B(n6032), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n59 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n101 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U61  ( .A(
        n8416), .B(n8871), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n58 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U60  ( .A(
        n8416), .B(n6032), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n58 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n100 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U59  ( .A(
        n8119), .B(n8871), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n57 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U58  ( .A(
        n8119), .B(n6032), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n57 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n99 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U57  ( .A(
        n7869), .B(n8871), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n56 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U56  ( .A(
        n7869), .B(n6032), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n56 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n98 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U55  ( .A(
        n7448), .B(n8871), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n54 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U54  ( .A(
        n7448), .B(n6032), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n54 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n97 ) );
  NAND3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U53  ( .A(
        recentABools_data_address0[3]), .B(recentABools_data_address0[4]), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n19 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n37 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U50  ( .A(
        n8870), .B(n7444), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n51 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U49  ( .A(
        n7653), .B(n7444), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n51 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n96 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U48  ( .A(
        n8870), .B(n6023), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n49 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U47  ( .A(
        n7653), .B(n6023), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n49 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n95 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U46  ( .A(
        n8870), .B(n6031), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n47 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U45  ( .A(
        n7653), .B(n6031), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n47 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n94 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U44  ( .A(
        n8870), .B(n6030), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n45 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U43  ( .A(
        n7653), .B(n6030), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n45 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n93 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U42  ( .A(
        n8870), .B(n8416), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n43 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U41  ( .A(
        n7653), .B(n8416), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n43 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n92 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U40  ( .A(
        n8870), .B(n8119), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n41 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U39  ( .A(
        n7653), .B(n8119), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n41 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n91 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U38  ( .A(
        n8870), .B(n7869), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n39 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U37  ( .A(
        n7653), .B(n7869), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n39 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n90 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U36  ( .A(
        n8870), .B(n7448), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n36 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U35  ( .A(
        n7448), .B(n7653), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n36 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n89 ) );
  AOI22X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U33  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n137 ), .B(
        recentABools_data_address0[2]), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n134 ), .D(n7648), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n30 ) );
  AOI22X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U32  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n131 ), .B(
        recentABools_data_address0[2]), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n128 ), .D(n7648), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n32 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U30  ( .A(
        n8402), .B(n6935), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n31 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n22 ) );
  AOI22X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U29  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n125 ), .B(
        recentABools_data_address0[2]), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n122 ), .D(n7648), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n25 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U27  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n140 ), .B(
        recentABools_data_address0[2]), .C(n6556), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n27 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U25  ( .A(
        n8402), .B(n7082), .C(n6555), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n24 ) );
  AOI22X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U24  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n22 ), .B(
        recentABools_data_address0[4]), .C(n6016), .D(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n24 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n21 ) );
  NOR3X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U23  ( .A(N461), 
        .B(ap_CS_fsm[9]), .C(n5902), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n20 ) );
  AOI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U22  ( .A(
        \tmp_12_reg_1694[0] ), .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n19 ), .C(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n20 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n16 ) );
  AOI22X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U18  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n159 ), .B(n8405), .C(\recentABools_data_U/Decision_recentVBools_data_ram_U/n156 ), .D(n10276), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n12 ) );
  AOI22X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U17  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n153 ), .B(n8405), .C(\recentABools_data_U/Decision_recentVBools_data_ram_U/n150 ), .D(n10276), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n15 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U14  ( .A(
        n10274), .B(n5696), .C(n4937), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n4 ) );
  AOI22X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U12  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n147 ), .B(n8405), .C(\recentABools_data_U/Decision_recentVBools_data_ram_U/n144 ), .D(n10276), 
        .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n7 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U10  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n162 ), .B(n8405), .C(n7967), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n9 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U8  ( .A(
        n10274), .B(n7594), .C(n7593), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n6 ) );
  AOI22X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U7  ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n4 ), .B(n7841), 
        .C(n10273), .D(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n6 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n1 ) );
  OAI21X1 \recentABools_data_U/Decision_recentVBools_data_ram_U/U4  ( .A(n7399), .B(n10534), .C(n7398), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n87 ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/q1_reg[0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n87 ), .CLK(
        n9069), .Q(\recentABools_data_q1[0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/q0_reg[0]  ( 
        .D(n4763), .CLK(n9069), .Q(\recentABools_data_q0[0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[0][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n89 ), .CLK(
        n9069), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[0][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[1][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n90 ), .CLK(
        n9069), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[1][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[2][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n91 ), .CLK(
        n9069), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[2][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[3][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n92 ), .CLK(
        n9069), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[3][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[4][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n93 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[4][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[5][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n94 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[5][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[6][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n95 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[6][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[7][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n96 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[7][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[8][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n97 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[8][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[9][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n98 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[9][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[10][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n99 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[10][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[11][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n100 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[11][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[12][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n101 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[12][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[13][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n102 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[13][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[14][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n103 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[14][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[15][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n104 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[15][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[16][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n105 ), .CLK(
        n9068), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[16][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[17][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n106 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[17][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[18][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n107 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[18][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[19][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n108 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[19][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[20][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n109 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[20][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[21][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n110 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[21][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[22][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n111 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[22][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[23][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n112 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[23][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[24][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n113 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[24][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[25][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n114 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[25][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[26][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n115 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[26][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[27][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n116 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[27][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[28][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n117 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[28][0] ) );
  DFFPOSX1 \recentABools_data_U/Decision_recentVBools_data_ram_U/ram_reg[29][0]  ( 
        .D(\recentABools_data_U/Decision_recentVBools_data_ram_U/n118 ), .CLK(
        n9067), .Q(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/ram[29][0] ) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_1  ( .A(\dp_cluster_1/N923 ), .B(
        \dp_cluster_1/N922 ), .YC(\dp_cluster_1/add_1107_aco/carry[2] ), .YS(
        tmp_6_fu_497_p3[1]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_2  ( .A(\dp_cluster_1/N924 ), .B(
        \dp_cluster_1/add_1107_aco/carry[2] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[3] ), .YS(tmp_6_fu_497_p3[2]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_3  ( .A(\dp_cluster_1/N925 ), .B(
        \dp_cluster_1/add_1107_aco/carry[3] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[4] ), .YS(tmp_6_fu_497_p3[3]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_4  ( .A(\dp_cluster_1/N926 ), .B(
        \dp_cluster_1/add_1107_aco/carry[4] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[5] ), .YS(tmp_6_fu_497_p3[4]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_5  ( .A(\dp_cluster_1/N927 ), .B(
        \dp_cluster_1/add_1107_aco/carry[5] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[6] ), .YS(tmp_6_fu_497_p3[5]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_6  ( .A(\dp_cluster_1/N928 ), .B(
        \dp_cluster_1/add_1107_aco/carry[6] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[7] ), .YS(tmp_6_fu_497_p3[6]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_7  ( .A(\dp_cluster_1/N929 ), .B(
        \dp_cluster_1/add_1107_aco/carry[7] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[8] ), .YS(tmp_6_fu_497_p3[7]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_8  ( .A(\dp_cluster_1/N930 ), .B(
        \dp_cluster_1/add_1107_aco/carry[8] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[9] ), .YS(tmp_6_fu_497_p3[8]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_9  ( .A(\dp_cluster_1/N931 ), .B(
        \dp_cluster_1/add_1107_aco/carry[9] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[10] ), .YS(tmp_6_fu_497_p3[9]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_10  ( .A(\dp_cluster_1/N932 ), .B(
        \dp_cluster_1/add_1107_aco/carry[10] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[11] ), .YS(tmp_6_fu_497_p3[10]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_11  ( .A(\dp_cluster_1/N933 ), .B(
        \dp_cluster_1/add_1107_aco/carry[11] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[12] ), .YS(tmp_6_fu_497_p3[11]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_12  ( .A(\dp_cluster_1/N934 ), .B(
        \dp_cluster_1/add_1107_aco/carry[12] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[13] ), .YS(tmp_6_fu_497_p3[12]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_13  ( .A(\dp_cluster_1/N935 ), .B(
        \dp_cluster_1/add_1107_aco/carry[13] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[14] ), .YS(tmp_6_fu_497_p3[13]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_14  ( .A(\dp_cluster_1/N936 ), .B(
        \dp_cluster_1/add_1107_aco/carry[14] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[15] ), .YS(tmp_6_fu_497_p3[14]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_15  ( .A(\dp_cluster_1/N937 ), .B(
        \dp_cluster_1/add_1107_aco/carry[15] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[16] ), .YS(tmp_6_fu_497_p3[15]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_16  ( .A(\dp_cluster_1/N938 ), .B(
        \dp_cluster_1/add_1107_aco/carry[16] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[17] ), .YS(tmp_6_fu_497_p3[16]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_17  ( .A(\dp_cluster_1/N939 ), .B(
        \dp_cluster_1/add_1107_aco/carry[17] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[18] ), .YS(tmp_6_fu_497_p3[17]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_18  ( .A(\dp_cluster_1/N940 ), .B(
        \dp_cluster_1/add_1107_aco/carry[18] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[19] ), .YS(tmp_6_fu_497_p3[18]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_19  ( .A(\dp_cluster_1/N941 ), .B(
        \dp_cluster_1/add_1107_aco/carry[19] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[20] ), .YS(tmp_6_fu_497_p3[19]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_20  ( .A(\dp_cluster_1/N942 ), .B(
        \dp_cluster_1/add_1107_aco/carry[20] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[21] ), .YS(tmp_6_fu_497_p3[20]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_21  ( .A(\dp_cluster_1/N943 ), .B(
        \dp_cluster_1/add_1107_aco/carry[21] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[22] ), .YS(tmp_6_fu_497_p3[21]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_22  ( .A(\dp_cluster_1/N944 ), .B(
        \dp_cluster_1/add_1107_aco/carry[22] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[23] ), .YS(tmp_6_fu_497_p3[22]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_23  ( .A(\dp_cluster_1/N945 ), .B(
        \dp_cluster_1/add_1107_aco/carry[23] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[24] ), .YS(tmp_6_fu_497_p3[23]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_24  ( .A(\dp_cluster_1/N946 ), .B(
        \dp_cluster_1/add_1107_aco/carry[24] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[25] ), .YS(tmp_6_fu_497_p3[24]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_25  ( .A(\dp_cluster_1/N947 ), .B(
        \dp_cluster_1/add_1107_aco/carry[25] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[26] ), .YS(tmp_6_fu_497_p3[25]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_26  ( .A(\dp_cluster_1/N948 ), .B(
        \dp_cluster_1/add_1107_aco/carry[26] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[27] ), .YS(tmp_6_fu_497_p3[26]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_27  ( .A(\dp_cluster_1/N949 ), .B(
        \dp_cluster_1/add_1107_aco/carry[27] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[28] ), .YS(tmp_6_fu_497_p3[27]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_28  ( .A(\dp_cluster_1/N950 ), .B(
        \dp_cluster_1/add_1107_aco/carry[28] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[29] ), .YS(tmp_6_fu_497_p3[28]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_29  ( .A(\dp_cluster_1/N951 ), .B(
        \dp_cluster_1/add_1107_aco/carry[29] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[30] ), .YS(tmp_6_fu_497_p3[29]) );
  HAX1 \dp_cluster_1/add_1107_aco/U1_1_30  ( .A(\dp_cluster_1/N952 ), .B(
        \dp_cluster_1/add_1107_aco/carry[30] ), .YC(
        \dp_cluster_1/add_1107_aco/carry[31] ), .YS(tmp_6_fu_497_p3[30]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_1  ( .A(\dp_cluster_0/N955 ), .B(
        \dp_cluster_0/N954 ), .YC(\dp_cluster_0/add_1147_aco/carry[2] ), .YS(
        tmp_7_fu_511_p3[1]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_2  ( .A(\dp_cluster_0/N956 ), .B(
        \dp_cluster_0/add_1147_aco/carry[2] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[3] ), .YS(tmp_7_fu_511_p3[2]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_3  ( .A(\dp_cluster_0/N957 ), .B(
        \dp_cluster_0/add_1147_aco/carry[3] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[4] ), .YS(tmp_7_fu_511_p3[3]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_4  ( .A(\dp_cluster_0/N958 ), .B(
        \dp_cluster_0/add_1147_aco/carry[4] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[5] ), .YS(tmp_7_fu_511_p3[4]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_5  ( .A(\dp_cluster_0/N959 ), .B(
        \dp_cluster_0/add_1147_aco/carry[5] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[6] ), .YS(tmp_7_fu_511_p3[5]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_6  ( .A(\dp_cluster_0/N960 ), .B(
        \dp_cluster_0/add_1147_aco/carry[6] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[7] ), .YS(tmp_7_fu_511_p3[6]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_7  ( .A(\dp_cluster_0/N961 ), .B(
        \dp_cluster_0/add_1147_aco/carry[7] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[8] ), .YS(tmp_7_fu_511_p3[7]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_8  ( .A(\dp_cluster_0/N962 ), .B(
        \dp_cluster_0/add_1147_aco/carry[8] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[9] ), .YS(tmp_7_fu_511_p3[8]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_9  ( .A(\dp_cluster_0/N963 ), .B(
        \dp_cluster_0/add_1147_aco/carry[9] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[10] ), .YS(tmp_7_fu_511_p3[9]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_10  ( .A(\dp_cluster_0/N964 ), .B(
        \dp_cluster_0/add_1147_aco/carry[10] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[11] ), .YS(tmp_7_fu_511_p3[10]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_11  ( .A(\dp_cluster_0/N965 ), .B(
        \dp_cluster_0/add_1147_aco/carry[11] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[12] ), .YS(tmp_7_fu_511_p3[11]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_12  ( .A(\dp_cluster_0/N966 ), .B(
        \dp_cluster_0/add_1147_aco/carry[12] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[13] ), .YS(tmp_7_fu_511_p3[12]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_13  ( .A(\dp_cluster_0/N967 ), .B(
        \dp_cluster_0/add_1147_aco/carry[13] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[14] ), .YS(tmp_7_fu_511_p3[13]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_14  ( .A(\dp_cluster_0/N968 ), .B(
        \dp_cluster_0/add_1147_aco/carry[14] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[15] ), .YS(tmp_7_fu_511_p3[14]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_15  ( .A(\dp_cluster_0/N969 ), .B(
        \dp_cluster_0/add_1147_aco/carry[15] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[16] ), .YS(tmp_7_fu_511_p3[15]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_16  ( .A(\dp_cluster_0/N970 ), .B(
        \dp_cluster_0/add_1147_aco/carry[16] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[17] ), .YS(tmp_7_fu_511_p3[16]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_17  ( .A(\dp_cluster_0/N971 ), .B(
        \dp_cluster_0/add_1147_aco/carry[17] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[18] ), .YS(tmp_7_fu_511_p3[17]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_18  ( .A(\dp_cluster_0/N972 ), .B(
        \dp_cluster_0/add_1147_aco/carry[18] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[19] ), .YS(tmp_7_fu_511_p3[18]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_19  ( .A(\dp_cluster_0/N973 ), .B(
        \dp_cluster_0/add_1147_aco/carry[19] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[20] ), .YS(tmp_7_fu_511_p3[19]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_20  ( .A(\dp_cluster_0/N974 ), .B(
        \dp_cluster_0/add_1147_aco/carry[20] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[21] ), .YS(tmp_7_fu_511_p3[20]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_21  ( .A(\dp_cluster_0/N975 ), .B(
        \dp_cluster_0/add_1147_aco/carry[21] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[22] ), .YS(tmp_7_fu_511_p3[21]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_22  ( .A(\dp_cluster_0/N976 ), .B(
        \dp_cluster_0/add_1147_aco/carry[22] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[23] ), .YS(tmp_7_fu_511_p3[22]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_23  ( .A(\dp_cluster_0/N977 ), .B(
        \dp_cluster_0/add_1147_aco/carry[23] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[24] ), .YS(tmp_7_fu_511_p3[23]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_24  ( .A(\dp_cluster_0/N978 ), .B(
        \dp_cluster_0/add_1147_aco/carry[24] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[25] ), .YS(tmp_7_fu_511_p3[24]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_25  ( .A(\dp_cluster_0/N979 ), .B(
        \dp_cluster_0/add_1147_aco/carry[25] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[26] ), .YS(tmp_7_fu_511_p3[25]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_26  ( .A(\dp_cluster_0/N980 ), .B(
        \dp_cluster_0/add_1147_aco/carry[26] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[27] ), .YS(tmp_7_fu_511_p3[26]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_27  ( .A(\dp_cluster_0/N981 ), .B(
        \dp_cluster_0/add_1147_aco/carry[27] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[28] ), .YS(tmp_7_fu_511_p3[27]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_28  ( .A(\dp_cluster_0/N982 ), .B(
        \dp_cluster_0/add_1147_aco/carry[28] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[29] ), .YS(tmp_7_fu_511_p3[28]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_29  ( .A(\dp_cluster_0/N983 ), .B(
        \dp_cluster_0/add_1147_aco/carry[29] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[30] ), .YS(tmp_7_fu_511_p3[29]) );
  HAX1 \dp_cluster_0/add_1147_aco/U1_1_30  ( .A(\dp_cluster_0/N984 ), .B(
        \dp_cluster_0/add_1147_aco/carry[30] ), .YC(
        \dp_cluster_0/add_1147_aco/carry[31] ), .YS(tmp_7_fu_511_p3[30]) );
  HAX1 \add_1415/U1_1_1  ( .A(VbeatFallDelay[1]), .B(VbeatFallDelay[0]), .YC(
        \add_1415/carry[2] ), .YS(tmp_5_fu_726_p2[1]) );
  HAX1 \add_1415/U1_1_2  ( .A(VbeatFallDelay[2]), .B(\add_1415/carry[2] ), 
        .YC(\add_1415/carry[3] ), .YS(tmp_5_fu_726_p2[2]) );
  HAX1 \add_1415/U1_1_3  ( .A(VbeatFallDelay[3]), .B(\add_1415/carry[3] ), 
        .YC(\add_1415/carry[4] ), .YS(tmp_5_fu_726_p2[3]) );
  HAX1 \add_1415/U1_1_4  ( .A(VbeatFallDelay[4]), .B(\add_1415/carry[4] ), 
        .YC(\add_1415/carry[5] ), .YS(tmp_5_fu_726_p2[4]) );
  HAX1 \add_1415/U1_1_5  ( .A(VbeatFallDelay[5]), .B(\add_1415/carry[5] ), 
        .YC(\add_1415/carry[6] ), .YS(tmp_5_fu_726_p2[5]) );
  HAX1 \add_1415/U1_1_6  ( .A(VbeatFallDelay[6]), .B(\add_1415/carry[6] ), 
        .YC(\add_1415/carry[7] ), .YS(tmp_5_fu_726_p2[6]) );
  HAX1 \add_1415/U1_1_7  ( .A(VbeatFallDelay[7]), .B(\add_1415/carry[7] ), 
        .YC(\add_1415/carry[8] ), .YS(tmp_5_fu_726_p2[7]) );
  HAX1 \add_1415/U1_1_8  ( .A(VbeatFallDelay[8]), .B(\add_1415/carry[8] ), 
        .YC(\add_1415/carry[9] ), .YS(tmp_5_fu_726_p2[8]) );
  HAX1 \add_1415/U1_1_9  ( .A(VbeatFallDelay[9]), .B(\add_1415/carry[9] ), 
        .YC(\add_1415/carry[10] ), .YS(tmp_5_fu_726_p2[9]) );
  HAX1 \add_1415/U1_1_10  ( .A(VbeatFallDelay[10]), .B(\add_1415/carry[10] ), 
        .YC(\add_1415/carry[11] ), .YS(tmp_5_fu_726_p2[10]) );
  HAX1 \add_1415/U1_1_11  ( .A(VbeatFallDelay[11]), .B(\add_1415/carry[11] ), 
        .YC(\add_1415/carry[12] ), .YS(tmp_5_fu_726_p2[11]) );
  HAX1 \add_1415/U1_1_12  ( .A(VbeatFallDelay[12]), .B(\add_1415/carry[12] ), 
        .YC(\add_1415/carry[13] ), .YS(tmp_5_fu_726_p2[12]) );
  HAX1 \add_1415/U1_1_13  ( .A(VbeatFallDelay[13]), .B(\add_1415/carry[13] ), 
        .YC(\add_1415/carry[14] ), .YS(tmp_5_fu_726_p2[13]) );
  HAX1 \add_1415/U1_1_14  ( .A(VbeatFallDelay[14]), .B(\add_1415/carry[14] ), 
        .YC(\add_1415/carry[15] ), .YS(tmp_5_fu_726_p2[14]) );
  HAX1 \add_1415/U1_1_15  ( .A(VbeatFallDelay[15]), .B(\add_1415/carry[15] ), 
        .YC(\add_1415/carry[16] ), .YS(tmp_5_fu_726_p2[15]) );
  HAX1 \add_1415/U1_1_16  ( .A(VbeatFallDelay[16]), .B(\add_1415/carry[16] ), 
        .YC(\add_1415/carry[17] ), .YS(tmp_5_fu_726_p2[16]) );
  HAX1 \add_1415/U1_1_17  ( .A(VbeatFallDelay[17]), .B(\add_1415/carry[17] ), 
        .YC(\add_1415/carry[18] ), .YS(tmp_5_fu_726_p2[17]) );
  HAX1 \add_1415/U1_1_18  ( .A(VbeatFallDelay[18]), .B(\add_1415/carry[18] ), 
        .YC(\add_1415/carry[19] ), .YS(tmp_5_fu_726_p2[18]) );
  HAX1 \add_1415/U1_1_19  ( .A(VbeatFallDelay[19]), .B(\add_1415/carry[19] ), 
        .YC(\add_1415/carry[20] ), .YS(tmp_5_fu_726_p2[19]) );
  HAX1 \add_1415/U1_1_20  ( .A(VbeatFallDelay[20]), .B(\add_1415/carry[20] ), 
        .YC(\add_1415/carry[21] ), .YS(tmp_5_fu_726_p2[20]) );
  HAX1 \add_1415/U1_1_21  ( .A(VbeatFallDelay[21]), .B(\add_1415/carry[21] ), 
        .YC(\add_1415/carry[22] ), .YS(tmp_5_fu_726_p2[21]) );
  HAX1 \add_1415/U1_1_22  ( .A(VbeatFallDelay[22]), .B(\add_1415/carry[22] ), 
        .YC(\add_1415/carry[23] ), .YS(tmp_5_fu_726_p2[22]) );
  HAX1 \add_1415/U1_1_23  ( .A(VbeatFallDelay[23]), .B(\add_1415/carry[23] ), 
        .YC(\add_1415/carry[24] ), .YS(tmp_5_fu_726_p2[23]) );
  HAX1 \add_1415/U1_1_24  ( .A(VbeatFallDelay[24]), .B(\add_1415/carry[24] ), 
        .YC(\add_1415/carry[25] ), .YS(tmp_5_fu_726_p2[24]) );
  HAX1 \add_1415/U1_1_25  ( .A(VbeatFallDelay[25]), .B(\add_1415/carry[25] ), 
        .YC(\add_1415/carry[26] ), .YS(tmp_5_fu_726_p2[25]) );
  HAX1 \add_1415/U1_1_26  ( .A(VbeatFallDelay[26]), .B(\add_1415/carry[26] ), 
        .YC(\add_1415/carry[27] ), .YS(tmp_5_fu_726_p2[26]) );
  HAX1 \add_1415/U1_1_27  ( .A(VbeatFallDelay[27]), .B(\add_1415/carry[27] ), 
        .YC(\add_1415/carry[28] ), .YS(tmp_5_fu_726_p2[27]) );
  HAX1 \add_1415/U1_1_28  ( .A(VbeatFallDelay[28]), .B(\add_1415/carry[28] ), 
        .YC(\add_1415/carry[29] ), .YS(tmp_5_fu_726_p2[28]) );
  HAX1 \add_1415/U1_1_29  ( .A(VbeatFallDelay[29]), .B(\add_1415/carry[29] ), 
        .YC(\add_1415/carry[30] ), .YS(tmp_5_fu_726_p2[29]) );
  HAX1 \add_1415/U1_1_30  ( .A(VbeatFallDelay[30]), .B(\add_1415/carry[30] ), 
        .YC(\add_1415/carry[31] ), .YS(tmp_5_fu_726_p2[30]) );
  HAX1 \add_1413/U1_1_1  ( .A(VbeatDelay[1]), .B(VbeatDelay[0]), .YC(
        \add_1413/carry[2] ), .YS(tmp_4_fu_716_p2[1]) );
  HAX1 \add_1413/U1_1_2  ( .A(VbeatDelay[2]), .B(\add_1413/carry[2] ), .YC(
        \add_1413/carry[3] ), .YS(tmp_4_fu_716_p2[2]) );
  HAX1 \add_1413/U1_1_3  ( .A(VbeatDelay[3]), .B(\add_1413/carry[3] ), .YC(
        \add_1413/carry[4] ), .YS(tmp_4_fu_716_p2[3]) );
  HAX1 \add_1413/U1_1_4  ( .A(VbeatDelay[4]), .B(\add_1413/carry[4] ), .YC(
        \add_1413/carry[5] ), .YS(tmp_4_fu_716_p2[4]) );
  HAX1 \add_1413/U1_1_5  ( .A(VbeatDelay[5]), .B(\add_1413/carry[5] ), .YC(
        \add_1413/carry[6] ), .YS(tmp_4_fu_716_p2[5]) );
  HAX1 \add_1413/U1_1_6  ( .A(VbeatDelay[6]), .B(\add_1413/carry[6] ), .YC(
        \add_1413/carry[7] ), .YS(tmp_4_fu_716_p2[6]) );
  HAX1 \add_1413/U1_1_7  ( .A(VbeatDelay[7]), .B(\add_1413/carry[7] ), .YC(
        \add_1413/carry[8] ), .YS(tmp_4_fu_716_p2[7]) );
  HAX1 \add_1413/U1_1_8  ( .A(VbeatDelay[8]), .B(\add_1413/carry[8] ), .YC(
        \add_1413/carry[9] ), .YS(tmp_4_fu_716_p2[8]) );
  HAX1 \add_1413/U1_1_9  ( .A(VbeatDelay[9]), .B(\add_1413/carry[9] ), .YC(
        \add_1413/carry[10] ), .YS(tmp_4_fu_716_p2[9]) );
  HAX1 \add_1413/U1_1_10  ( .A(VbeatDelay[10]), .B(\add_1413/carry[10] ), .YC(
        \add_1413/carry[11] ), .YS(tmp_4_fu_716_p2[10]) );
  HAX1 \add_1413/U1_1_11  ( .A(VbeatDelay[11]), .B(\add_1413/carry[11] ), .YC(
        \add_1413/carry[12] ), .YS(tmp_4_fu_716_p2[11]) );
  HAX1 \add_1413/U1_1_12  ( .A(VbeatDelay[12]), .B(\add_1413/carry[12] ), .YC(
        \add_1413/carry[13] ), .YS(tmp_4_fu_716_p2[12]) );
  HAX1 \add_1413/U1_1_13  ( .A(VbeatDelay[13]), .B(\add_1413/carry[13] ), .YC(
        \add_1413/carry[14] ), .YS(tmp_4_fu_716_p2[13]) );
  HAX1 \add_1413/U1_1_14  ( .A(VbeatDelay[14]), .B(\add_1413/carry[14] ), .YC(
        \add_1413/carry[15] ), .YS(tmp_4_fu_716_p2[14]) );
  HAX1 \add_1413/U1_1_15  ( .A(VbeatDelay[15]), .B(\add_1413/carry[15] ), .YC(
        \add_1413/carry[16] ), .YS(tmp_4_fu_716_p2[15]) );
  HAX1 \add_1413/U1_1_16  ( .A(VbeatDelay[16]), .B(\add_1413/carry[16] ), .YC(
        \add_1413/carry[17] ), .YS(tmp_4_fu_716_p2[16]) );
  HAX1 \add_1413/U1_1_17  ( .A(VbeatDelay[17]), .B(\add_1413/carry[17] ), .YC(
        \add_1413/carry[18] ), .YS(tmp_4_fu_716_p2[17]) );
  HAX1 \add_1413/U1_1_18  ( .A(VbeatDelay[18]), .B(\add_1413/carry[18] ), .YC(
        \add_1413/carry[19] ), .YS(tmp_4_fu_716_p2[18]) );
  HAX1 \add_1413/U1_1_19  ( .A(VbeatDelay[19]), .B(\add_1413/carry[19] ), .YC(
        \add_1413/carry[20] ), .YS(tmp_4_fu_716_p2[19]) );
  HAX1 \add_1413/U1_1_20  ( .A(VbeatDelay[20]), .B(\add_1413/carry[20] ), .YC(
        \add_1413/carry[21] ), .YS(tmp_4_fu_716_p2[20]) );
  HAX1 \add_1413/U1_1_21  ( .A(VbeatDelay[21]), .B(\add_1413/carry[21] ), .YC(
        \add_1413/carry[22] ), .YS(tmp_4_fu_716_p2[21]) );
  HAX1 \add_1413/U1_1_22  ( .A(VbeatDelay[22]), .B(\add_1413/carry[22] ), .YC(
        \add_1413/carry[23] ), .YS(tmp_4_fu_716_p2[22]) );
  HAX1 \add_1413/U1_1_23  ( .A(VbeatDelay[23]), .B(\add_1413/carry[23] ), .YC(
        \add_1413/carry[24] ), .YS(tmp_4_fu_716_p2[23]) );
  HAX1 \add_1413/U1_1_24  ( .A(VbeatDelay[24]), .B(\add_1413/carry[24] ), .YC(
        \add_1413/carry[25] ), .YS(tmp_4_fu_716_p2[24]) );
  HAX1 \add_1413/U1_1_25  ( .A(VbeatDelay[25]), .B(\add_1413/carry[25] ), .YC(
        \add_1413/carry[26] ), .YS(tmp_4_fu_716_p2[25]) );
  HAX1 \add_1413/U1_1_26  ( .A(VbeatDelay[26]), .B(\add_1413/carry[26] ), .YC(
        \add_1413/carry[27] ), .YS(tmp_4_fu_716_p2[26]) );
  HAX1 \add_1413/U1_1_27  ( .A(VbeatDelay[27]), .B(\add_1413/carry[27] ), .YC(
        \add_1413/carry[28] ), .YS(tmp_4_fu_716_p2[27]) );
  HAX1 \add_1413/U1_1_28  ( .A(VbeatDelay[28]), .B(\add_1413/carry[28] ), .YC(
        \add_1413/carry[29] ), .YS(tmp_4_fu_716_p2[28]) );
  HAX1 \add_1413/U1_1_29  ( .A(VbeatDelay[29]), .B(\add_1413/carry[29] ), .YC(
        \add_1413/carry[30] ), .YS(tmp_4_fu_716_p2[29]) );
  HAX1 \add_1413/U1_1_30  ( .A(VbeatDelay[30]), .B(\add_1413/carry[30] ), .YC(
        \add_1413/carry[31] ), .YS(tmp_4_fu_716_p2[30]) );
  HAX1 \add_1407/U1_1_1  ( .A(AbeatDelay[1]), .B(AbeatDelay[0]), .YC(
        \add_1407/carry[2] ), .YS(tmp_3_fu_706_p2[1]) );
  HAX1 \add_1407/U1_1_2  ( .A(AbeatDelay[2]), .B(\add_1407/carry[2] ), .YC(
        \add_1407/carry[3] ), .YS(tmp_3_fu_706_p2[2]) );
  HAX1 \add_1407/U1_1_3  ( .A(AbeatDelay[3]), .B(\add_1407/carry[3] ), .YC(
        \add_1407/carry[4] ), .YS(tmp_3_fu_706_p2[3]) );
  HAX1 \add_1407/U1_1_4  ( .A(AbeatDelay[4]), .B(\add_1407/carry[4] ), .YC(
        \add_1407/carry[5] ), .YS(tmp_3_fu_706_p2[4]) );
  HAX1 \add_1407/U1_1_5  ( .A(AbeatDelay[5]), .B(\add_1407/carry[5] ), .YC(
        \add_1407/carry[6] ), .YS(tmp_3_fu_706_p2[5]) );
  HAX1 \add_1407/U1_1_6  ( .A(AbeatDelay[6]), .B(\add_1407/carry[6] ), .YC(
        \add_1407/carry[7] ), .YS(tmp_3_fu_706_p2[6]) );
  HAX1 \add_1407/U1_1_7  ( .A(AbeatDelay[7]), .B(\add_1407/carry[7] ), .YC(
        \add_1407/carry[8] ), .YS(tmp_3_fu_706_p2[7]) );
  HAX1 \add_1407/U1_1_8  ( .A(AbeatDelay[8]), .B(\add_1407/carry[8] ), .YC(
        \add_1407/carry[9] ), .YS(tmp_3_fu_706_p2[8]) );
  HAX1 \add_1407/U1_1_9  ( .A(AbeatDelay[9]), .B(\add_1407/carry[9] ), .YC(
        \add_1407/carry[10] ), .YS(tmp_3_fu_706_p2[9]) );
  HAX1 \add_1407/U1_1_10  ( .A(AbeatDelay[10]), .B(\add_1407/carry[10] ), .YC(
        \add_1407/carry[11] ), .YS(tmp_3_fu_706_p2[10]) );
  HAX1 \add_1407/U1_1_11  ( .A(AbeatDelay[11]), .B(\add_1407/carry[11] ), .YC(
        \add_1407/carry[12] ), .YS(tmp_3_fu_706_p2[11]) );
  HAX1 \add_1407/U1_1_12  ( .A(AbeatDelay[12]), .B(\add_1407/carry[12] ), .YC(
        \add_1407/carry[13] ), .YS(tmp_3_fu_706_p2[12]) );
  HAX1 \add_1407/U1_1_13  ( .A(AbeatDelay[13]), .B(\add_1407/carry[13] ), .YC(
        \add_1407/carry[14] ), .YS(tmp_3_fu_706_p2[13]) );
  HAX1 \add_1407/U1_1_14  ( .A(AbeatDelay[14]), .B(\add_1407/carry[14] ), .YC(
        \add_1407/carry[15] ), .YS(tmp_3_fu_706_p2[14]) );
  HAX1 \add_1407/U1_1_15  ( .A(AbeatDelay[15]), .B(\add_1407/carry[15] ), .YC(
        \add_1407/carry[16] ), .YS(tmp_3_fu_706_p2[15]) );
  HAX1 \add_1407/U1_1_16  ( .A(AbeatDelay[16]), .B(\add_1407/carry[16] ), .YC(
        \add_1407/carry[17] ), .YS(tmp_3_fu_706_p2[16]) );
  HAX1 \add_1407/U1_1_17  ( .A(AbeatDelay[17]), .B(\add_1407/carry[17] ), .YC(
        \add_1407/carry[18] ), .YS(tmp_3_fu_706_p2[17]) );
  HAX1 \add_1407/U1_1_18  ( .A(AbeatDelay[18]), .B(\add_1407/carry[18] ), .YC(
        \add_1407/carry[19] ), .YS(tmp_3_fu_706_p2[18]) );
  HAX1 \add_1407/U1_1_19  ( .A(AbeatDelay[19]), .B(\add_1407/carry[19] ), .YC(
        \add_1407/carry[20] ), .YS(tmp_3_fu_706_p2[19]) );
  HAX1 \add_1407/U1_1_20  ( .A(AbeatDelay[20]), .B(\add_1407/carry[20] ), .YC(
        \add_1407/carry[21] ), .YS(tmp_3_fu_706_p2[20]) );
  HAX1 \add_1407/U1_1_21  ( .A(AbeatDelay[21]), .B(\add_1407/carry[21] ), .YC(
        \add_1407/carry[22] ), .YS(tmp_3_fu_706_p2[21]) );
  HAX1 \add_1407/U1_1_22  ( .A(AbeatDelay[22]), .B(\add_1407/carry[22] ), .YC(
        \add_1407/carry[23] ), .YS(tmp_3_fu_706_p2[22]) );
  HAX1 \add_1407/U1_1_23  ( .A(AbeatDelay[23]), .B(\add_1407/carry[23] ), .YC(
        \add_1407/carry[24] ), .YS(tmp_3_fu_706_p2[23]) );
  HAX1 \add_1407/U1_1_24  ( .A(AbeatDelay[24]), .B(\add_1407/carry[24] ), .YC(
        \add_1407/carry[25] ), .YS(tmp_3_fu_706_p2[24]) );
  HAX1 \add_1407/U1_1_25  ( .A(AbeatDelay[25]), .B(\add_1407/carry[25] ), .YC(
        \add_1407/carry[26] ), .YS(tmp_3_fu_706_p2[25]) );
  HAX1 \add_1407/U1_1_26  ( .A(AbeatDelay[26]), .B(\add_1407/carry[26] ), .YC(
        \add_1407/carry[27] ), .YS(tmp_3_fu_706_p2[26]) );
  HAX1 \add_1407/U1_1_27  ( .A(AbeatDelay[27]), .B(\add_1407/carry[27] ), .YC(
        \add_1407/carry[28] ), .YS(tmp_3_fu_706_p2[27]) );
  HAX1 \add_1407/U1_1_28  ( .A(AbeatDelay[28]), .B(\add_1407/carry[28] ), .YC(
        \add_1407/carry[29] ), .YS(tmp_3_fu_706_p2[28]) );
  HAX1 \add_1407/U1_1_29  ( .A(AbeatDelay[29]), .B(\add_1407/carry[29] ), .YC(
        \add_1407/carry[30] ), .YS(tmp_3_fu_706_p2[29]) );
  HAX1 \add_1407/U1_1_30  ( .A(AbeatDelay[30]), .B(\add_1407/carry[30] ), .YC(
        \add_1407/carry[31] ), .YS(tmp_3_fu_706_p2[30]) );
  HAX1 \add_1405/U1_1_1  ( .A(recentdatapoints_head_i[1]), .B(
        recentdatapoints_head_i[0]), .YC(\add_1405/carry[2] ), .YS(
        p_tmp_i_fu_587_p3[1]) );
  HAX1 \add_1405/U1_1_2  ( .A(recentdatapoints_head_i[2]), .B(
        \add_1405/carry[2] ), .YC(\add_1405/carry[3] ), .YS(
        tmp_39_i_fu_576_p2[2]) );
  HAX1 \add_1405/U1_1_3  ( .A(recentdatapoints_head_i[3]), .B(
        \add_1405/carry[3] ), .YC(\add_1405/carry[4] ), .YS(
        p_tmp_i_fu_587_p3[3]) );
  HAX1 \add_1405/U1_1_4  ( .A(recentdatapoints_head_i[4]), .B(
        \add_1405/carry[4] ), .YC(\add_1405/carry[5] ), .YS(
        tmp_39_i_fu_576_p2[4]) );
  HAX1 \add_1405/U1_1_5  ( .A(recentdatapoints_head_i[5]), .B(
        \add_1405/carry[5] ), .YC(\add_1405/carry[6] ), .YS(
        p_tmp_i_fu_587_p3[5]) );
  HAX1 \add_1405/U1_1_6  ( .A(recentdatapoints_head_i[6]), .B(
        \add_1405/carry[6] ), .YC(\add_1405/carry[7] ), .YS(
        p_tmp_i_fu_587_p3[6]) );
  HAX1 \add_1405/U1_1_7  ( .A(recentdatapoints_head_i[7]), .B(
        \add_1405/carry[7] ), .YC(\add_1405/carry[8] ), .YS(
        p_tmp_i_fu_587_p3[7]) );
  HAX1 \add_1405/U1_1_8  ( .A(recentdatapoints_head_i[8]), .B(
        \add_1405/carry[8] ), .YC(\add_1405/carry[9] ), .YS(
        p_tmp_i_fu_587_p3[8]) );
  HAX1 \add_1405/U1_1_9  ( .A(recentdatapoints_head_i[9]), .B(
        \add_1405/carry[9] ), .YC(\add_1405/carry[10] ), .YS(
        p_tmp_i_fu_587_p3[9]) );
  HAX1 \add_1405/U1_1_10  ( .A(recentdatapoints_head_i[10]), .B(
        \add_1405/carry[10] ), .YC(\add_1405/carry[11] ), .YS(
        p_tmp_i_fu_587_p3[10]) );
  HAX1 \add_1405/U1_1_11  ( .A(recentdatapoints_head_i[11]), .B(
        \add_1405/carry[11] ), .YC(\add_1405/carry[12] ), .YS(
        p_tmp_i_fu_587_p3[11]) );
  HAX1 \add_1405/U1_1_12  ( .A(recentdatapoints_head_i[12]), .B(
        \add_1405/carry[12] ), .YC(\add_1405/carry[13] ), .YS(
        p_tmp_i_fu_587_p3[12]) );
  HAX1 \add_1405/U1_1_13  ( .A(recentdatapoints_head_i[13]), .B(
        \add_1405/carry[13] ), .YC(\add_1405/carry[14] ), .YS(
        p_tmp_i_fu_587_p3[13]) );
  HAX1 \add_1405/U1_1_14  ( .A(recentdatapoints_head_i[14]), .B(
        \add_1405/carry[14] ), .YC(\add_1405/carry[15] ), .YS(
        p_tmp_i_fu_587_p3[14]) );
  HAX1 \add_1405/U1_1_15  ( .A(recentdatapoints_head_i[15]), .B(
        \add_1405/carry[15] ), .YC(\add_1405/carry[16] ), .YS(
        p_tmp_i_fu_587_p3[15]) );
  HAX1 \add_1405/U1_1_16  ( .A(recentdatapoints_head_i[16]), .B(
        \add_1405/carry[16] ), .YC(\add_1405/carry[17] ), .YS(
        p_tmp_i_fu_587_p3[16]) );
  HAX1 \add_1405/U1_1_17  ( .A(recentdatapoints_head_i[17]), .B(
        \add_1405/carry[17] ), .YC(\add_1405/carry[18] ), .YS(
        p_tmp_i_fu_587_p3[17]) );
  HAX1 \add_1405/U1_1_18  ( .A(recentdatapoints_head_i[18]), .B(
        \add_1405/carry[18] ), .YC(\add_1405/carry[19] ), .YS(
        p_tmp_i_fu_587_p3[18]) );
  HAX1 \add_1405/U1_1_19  ( .A(recentdatapoints_head_i[19]), .B(
        \add_1405/carry[19] ), .YC(\add_1405/carry[20] ), .YS(
        p_tmp_i_fu_587_p3[19]) );
  HAX1 \add_1405/U1_1_20  ( .A(recentdatapoints_head_i[20]), .B(
        \add_1405/carry[20] ), .YC(\add_1405/carry[21] ), .YS(
        p_tmp_i_fu_587_p3[20]) );
  HAX1 \add_1405/U1_1_21  ( .A(recentdatapoints_head_i[21]), .B(
        \add_1405/carry[21] ), .YC(\add_1405/carry[22] ), .YS(
        p_tmp_i_fu_587_p3[21]) );
  HAX1 \add_1405/U1_1_22  ( .A(recentdatapoints_head_i[22]), .B(
        \add_1405/carry[22] ), .YC(\add_1405/carry[23] ), .YS(
        p_tmp_i_fu_587_p3[22]) );
  HAX1 \add_1405/U1_1_23  ( .A(recentdatapoints_head_i[23]), .B(
        \add_1405/carry[23] ), .YC(\add_1405/carry[24] ), .YS(
        p_tmp_i_fu_587_p3[23]) );
  HAX1 \add_1405/U1_1_24  ( .A(recentdatapoints_head_i[24]), .B(
        \add_1405/carry[24] ), .YC(\add_1405/carry[25] ), .YS(
        p_tmp_i_fu_587_p3[24]) );
  HAX1 \add_1405/U1_1_25  ( .A(recentdatapoints_head_i[25]), .B(
        \add_1405/carry[25] ), .YC(\add_1405/carry[26] ), .YS(
        p_tmp_i_fu_587_p3[25]) );
  HAX1 \add_1405/U1_1_26  ( .A(recentdatapoints_head_i[26]), .B(
        \add_1405/carry[26] ), .YC(\add_1405/carry[27] ), .YS(
        p_tmp_i_fu_587_p3[26]) );
  HAX1 \add_1405/U1_1_27  ( .A(recentdatapoints_head_i[27]), .B(
        \add_1405/carry[27] ), .YC(\add_1405/carry[28] ), .YS(
        p_tmp_i_fu_587_p3[27]) );
  HAX1 \add_1405/U1_1_28  ( .A(recentdatapoints_head_i[28]), .B(
        \add_1405/carry[28] ), .YC(\add_1405/carry[29] ), .YS(
        p_tmp_i_fu_587_p3[28]) );
  HAX1 \add_1405/U1_1_29  ( .A(recentdatapoints_head_i[29]), .B(
        \add_1405/carry[29] ), .YC(\add_1405/carry[30] ), .YS(
        p_tmp_i_fu_587_p3[29]) );
  HAX1 \add_1405/U1_1_30  ( .A(recentdatapoints_head_i[30]), .B(
        \add_1405/carry[30] ), .YC(\add_1405/carry[31] ), .YS(
        p_tmp_i_fu_587_p3[30]) );
  HAX1 \add_1393/U1_1_1  ( .A(recentVBools_head_i[1]), .B(
        recentVBools_head_i[0]), .YC(\add_1393/carry[2] ), .YS(
        tmp_33_i_fu_786_p2[1]) );
  HAX1 \add_1393/U1_1_2  ( .A(recentVBools_head_i[2]), .B(\add_1393/carry[2] ), 
        .YC(\add_1393/carry[3] ), .YS(tmp_33_i_fu_786_p2[2]) );
  HAX1 \add_1393/U1_1_3  ( .A(recentVBools_head_i[3]), .B(\add_1393/carry[3] ), 
        .YC(\add_1393/carry[4] ), .YS(tmp_33_i_fu_786_p2[3]) );
  HAX1 \add_1393/U1_1_4  ( .A(recentVBools_head_i[4]), .B(\add_1393/carry[4] ), 
        .YC(\add_1393/carry[5] ), .YS(tmp_33_i_fu_786_p2[4]) );
  HAX1 \add_1393/U1_1_5  ( .A(recentVBools_head_i[5]), .B(\add_1393/carry[5] ), 
        .YC(\add_1393/carry[6] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[5]) );
  HAX1 \add_1393/U1_1_6  ( .A(recentVBools_head_i[6]), .B(\add_1393/carry[6] ), 
        .YC(\add_1393/carry[7] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[6]) );
  HAX1 \add_1393/U1_1_7  ( .A(recentVBools_head_i[7]), .B(\add_1393/carry[7] ), 
        .YC(\add_1393/carry[8] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[7]) );
  HAX1 \add_1393/U1_1_8  ( .A(recentVBools_head_i[8]), .B(\add_1393/carry[8] ), 
        .YC(\add_1393/carry[9] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[8]) );
  HAX1 \add_1393/U1_1_9  ( .A(recentVBools_head_i[9]), .B(\add_1393/carry[9] ), 
        .YC(\add_1393/carry[10] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[9]) );
  HAX1 \add_1393/U1_1_10  ( .A(recentVBools_head_i[10]), .B(
        \add_1393/carry[10] ), .YC(\add_1393/carry[11] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[10]) );
  HAX1 \add_1393/U1_1_11  ( .A(recentVBools_head_i[11]), .B(
        \add_1393/carry[11] ), .YC(\add_1393/carry[12] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[11]) );
  HAX1 \add_1393/U1_1_12  ( .A(recentVBools_head_i[12]), .B(
        \add_1393/carry[12] ), .YC(\add_1393/carry[13] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[12]) );
  HAX1 \add_1393/U1_1_13  ( .A(recentVBools_head_i[13]), .B(
        \add_1393/carry[13] ), .YC(\add_1393/carry[14] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[13]) );
  HAX1 \add_1393/U1_1_14  ( .A(recentVBools_head_i[14]), .B(
        \add_1393/carry[14] ), .YC(\add_1393/carry[15] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[14]) );
  HAX1 \add_1393/U1_1_15  ( .A(recentVBools_head_i[15]), .B(
        \add_1393/carry[15] ), .YC(\add_1393/carry[16] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[15]) );
  HAX1 \add_1393/U1_1_16  ( .A(recentVBools_head_i[16]), .B(
        \add_1393/carry[16] ), .YC(\add_1393/carry[17] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[16]) );
  HAX1 \add_1393/U1_1_17  ( .A(recentVBools_head_i[17]), .B(
        \add_1393/carry[17] ), .YC(\add_1393/carry[18] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[17]) );
  HAX1 \add_1393/U1_1_18  ( .A(recentVBools_head_i[18]), .B(
        \add_1393/carry[18] ), .YC(\add_1393/carry[19] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[18]) );
  HAX1 \add_1393/U1_1_19  ( .A(recentVBools_head_i[19]), .B(
        \add_1393/carry[19] ), .YC(\add_1393/carry[20] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[19]) );
  HAX1 \add_1393/U1_1_20  ( .A(recentVBools_head_i[20]), .B(
        \add_1393/carry[20] ), .YC(\add_1393/carry[21] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[20]) );
  HAX1 \add_1393/U1_1_21  ( .A(recentVBools_head_i[21]), .B(
        \add_1393/carry[21] ), .YC(\add_1393/carry[22] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[21]) );
  HAX1 \add_1393/U1_1_22  ( .A(recentVBools_head_i[22]), .B(
        \add_1393/carry[22] ), .YC(\add_1393/carry[23] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[22]) );
  HAX1 \add_1393/U1_1_23  ( .A(recentVBools_head_i[23]), .B(
        \add_1393/carry[23] ), .YC(\add_1393/carry[24] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[23]) );
  HAX1 \add_1393/U1_1_24  ( .A(recentVBools_head_i[24]), .B(
        \add_1393/carry[24] ), .YC(\add_1393/carry[25] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[24]) );
  HAX1 \add_1393/U1_1_25  ( .A(recentVBools_head_i[25]), .B(
        \add_1393/carry[25] ), .YC(\add_1393/carry[26] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[25]) );
  HAX1 \add_1393/U1_1_26  ( .A(recentVBools_head_i[26]), .B(
        \add_1393/carry[26] ), .YC(\add_1393/carry[27] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[26]) );
  HAX1 \add_1393/U1_1_27  ( .A(recentVBools_head_i[27]), .B(
        \add_1393/carry[27] ), .YC(\add_1393/carry[28] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[27]) );
  HAX1 \add_1393/U1_1_28  ( .A(recentVBools_head_i[28]), .B(
        \add_1393/carry[28] ), .YC(\add_1393/carry[29] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[28]) );
  HAX1 \add_1393/U1_1_29  ( .A(recentVBools_head_i[29]), .B(
        \add_1393/carry[29] ), .YC(\add_1393/carry[30] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[29]) );
  HAX1 \add_1393/U1_1_30  ( .A(recentVBools_head_i[30]), .B(
        \add_1393/carry[30] ), .YC(\add_1393/carry[31] ), .YS(
        CircularBuffer_head_i_read_ass_fu_797_p3[30]) );
  HAX1 \add_1391/U1_1_1  ( .A(recentABools_head_i[1]), .B(
        recentABools_head_i[0]), .YC(\add_1391/carry[2] ), .YS(
        tmp_33_i1_fu_1099_p2[1]) );
  HAX1 \add_1391/U1_1_2  ( .A(recentABools_head_i[2]), .B(\add_1391/carry[2] ), 
        .YC(\add_1391/carry[3] ), .YS(tmp_33_i1_fu_1099_p2[2]) );
  HAX1 \add_1391/U1_1_3  ( .A(recentABools_head_i[3]), .B(\add_1391/carry[3] ), 
        .YC(\add_1391/carry[4] ), .YS(tmp_33_i1_fu_1099_p2[3]) );
  HAX1 \add_1391/U1_1_4  ( .A(recentABools_head_i[4]), .B(\add_1391/carry[4] ), 
        .YC(\add_1391/carry[5] ), .YS(tmp_33_i1_fu_1099_p2[4]) );
  HAX1 \add_1391/U1_1_5  ( .A(recentABools_head_i[5]), .B(\add_1391/carry[5] ), 
        .YC(\add_1391/carry[6] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[5]) );
  HAX1 \add_1391/U1_1_6  ( .A(recentABools_head_i[6]), .B(\add_1391/carry[6] ), 
        .YC(\add_1391/carry[7] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[6]) );
  HAX1 \add_1391/U1_1_7  ( .A(recentABools_head_i[7]), .B(\add_1391/carry[7] ), 
        .YC(\add_1391/carry[8] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[7]) );
  HAX1 \add_1391/U1_1_8  ( .A(recentABools_head_i[8]), .B(\add_1391/carry[8] ), 
        .YC(\add_1391/carry[9] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[8]) );
  HAX1 \add_1391/U1_1_9  ( .A(recentABools_head_i[9]), .B(\add_1391/carry[9] ), 
        .YC(\add_1391/carry[10] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[9]) );
  HAX1 \add_1391/U1_1_10  ( .A(recentABools_head_i[10]), .B(
        \add_1391/carry[10] ), .YC(\add_1391/carry[11] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[10]) );
  HAX1 \add_1391/U1_1_11  ( .A(recentABools_head_i[11]), .B(
        \add_1391/carry[11] ), .YC(\add_1391/carry[12] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[11]) );
  HAX1 \add_1391/U1_1_12  ( .A(recentABools_head_i[12]), .B(
        \add_1391/carry[12] ), .YC(\add_1391/carry[13] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[12]) );
  HAX1 \add_1391/U1_1_13  ( .A(recentABools_head_i[13]), .B(
        \add_1391/carry[13] ), .YC(\add_1391/carry[14] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[13]) );
  HAX1 \add_1391/U1_1_14  ( .A(recentABools_head_i[14]), .B(
        \add_1391/carry[14] ), .YC(\add_1391/carry[15] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[14]) );
  HAX1 \add_1391/U1_1_15  ( .A(recentABools_head_i[15]), .B(
        \add_1391/carry[15] ), .YC(\add_1391/carry[16] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[15]) );
  HAX1 \add_1391/U1_1_16  ( .A(recentABools_head_i[16]), .B(
        \add_1391/carry[16] ), .YC(\add_1391/carry[17] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[16]) );
  HAX1 \add_1391/U1_1_17  ( .A(recentABools_head_i[17]), .B(
        \add_1391/carry[17] ), .YC(\add_1391/carry[18] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[17]) );
  HAX1 \add_1391/U1_1_18  ( .A(recentABools_head_i[18]), .B(
        \add_1391/carry[18] ), .YC(\add_1391/carry[19] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[18]) );
  HAX1 \add_1391/U1_1_19  ( .A(recentABools_head_i[19]), .B(
        \add_1391/carry[19] ), .YC(\add_1391/carry[20] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[19]) );
  HAX1 \add_1391/U1_1_20  ( .A(recentABools_head_i[20]), .B(
        \add_1391/carry[20] ), .YC(\add_1391/carry[21] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[20]) );
  HAX1 \add_1391/U1_1_21  ( .A(recentABools_head_i[21]), .B(
        \add_1391/carry[21] ), .YC(\add_1391/carry[22] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[21]) );
  HAX1 \add_1391/U1_1_22  ( .A(recentABools_head_i[22]), .B(
        \add_1391/carry[22] ), .YC(\add_1391/carry[23] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[22]) );
  HAX1 \add_1391/U1_1_23  ( .A(recentABools_head_i[23]), .B(
        \add_1391/carry[23] ), .YC(\add_1391/carry[24] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[23]) );
  HAX1 \add_1391/U1_1_24  ( .A(recentABools_head_i[24]), .B(
        \add_1391/carry[24] ), .YC(\add_1391/carry[25] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[24]) );
  HAX1 \add_1391/U1_1_25  ( .A(recentABools_head_i[25]), .B(
        \add_1391/carry[25] ), .YC(\add_1391/carry[26] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[25]) );
  HAX1 \add_1391/U1_1_26  ( .A(recentABools_head_i[26]), .B(
        \add_1391/carry[26] ), .YC(\add_1391/carry[27] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[26]) );
  HAX1 \add_1391/U1_1_27  ( .A(recentABools_head_i[27]), .B(
        \add_1391/carry[27] ), .YC(\add_1391/carry[28] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[27]) );
  HAX1 \add_1391/U1_1_28  ( .A(recentABools_head_i[28]), .B(
        \add_1391/carry[28] ), .YC(\add_1391/carry[29] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[28]) );
  HAX1 \add_1391/U1_1_29  ( .A(recentABools_head_i[29]), .B(
        \add_1391/carry[29] ), .YC(\add_1391/carry[30] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[29]) );
  HAX1 \add_1391/U1_1_30  ( .A(recentABools_head_i[30]), .B(
        \add_1391/carry[30] ), .YC(\add_1391/carry[31] ), .YS(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[30]) );
  HAX1 \add_1319/U1_1_1  ( .A(recentdatapoints_len[1]), .B(
        recentdatapoints_len[0]), .YC(\add_1319/carry[2] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[1]) );
  HAX1 \add_1319/U1_1_2  ( .A(recentdatapoints_len[2]), .B(\add_1319/carry[2] ), .YC(\add_1319/carry[3] ), .YS(recentdatapoints_len_load_op_fu_556_p2[2]) );
  HAX1 \add_1319/U1_1_3  ( .A(recentdatapoints_len[3]), .B(\add_1319/carry[3] ), .YC(\add_1319/carry[4] ), .YS(recentdatapoints_len_load_op_fu_556_p2[3]) );
  HAX1 \add_1319/U1_1_4  ( .A(recentdatapoints_len[4]), .B(\add_1319/carry[4] ), .YC(\add_1319/carry[5] ), .YS(recentdatapoints_len_load_op_fu_556_p2[4]) );
  HAX1 \add_1319/U1_1_5  ( .A(recentdatapoints_len[5]), .B(\add_1319/carry[5] ), .YC(\add_1319/carry[6] ), .YS(recentdatapoints_len_load_op_fu_556_p2[5]) );
  HAX1 \add_1319/U1_1_6  ( .A(recentdatapoints_len[6]), .B(\add_1319/carry[6] ), .YC(\add_1319/carry[7] ), .YS(recentdatapoints_len_load_op_fu_556_p2[6]) );
  HAX1 \add_1319/U1_1_7  ( .A(recentdatapoints_len[7]), .B(\add_1319/carry[7] ), .YC(\add_1319/carry[8] ), .YS(recentdatapoints_len_load_op_fu_556_p2[7]) );
  HAX1 \add_1319/U1_1_8  ( .A(recentdatapoints_len[8]), .B(\add_1319/carry[8] ), .YC(\add_1319/carry[9] ), .YS(recentdatapoints_len_load_op_fu_556_p2[8]) );
  HAX1 \add_1319/U1_1_9  ( .A(recentdatapoints_len[9]), .B(\add_1319/carry[9] ), .YC(\add_1319/carry[10] ), .YS(recentdatapoints_len_load_op_fu_556_p2[9]) );
  HAX1 \add_1319/U1_1_10  ( .A(recentdatapoints_len[10]), .B(
        \add_1319/carry[10] ), .YC(\add_1319/carry[11] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[10]) );
  HAX1 \add_1319/U1_1_11  ( .A(recentdatapoints_len[11]), .B(
        \add_1319/carry[11] ), .YC(\add_1319/carry[12] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[11]) );
  HAX1 \add_1319/U1_1_12  ( .A(recentdatapoints_len[12]), .B(
        \add_1319/carry[12] ), .YC(\add_1319/carry[13] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[12]) );
  HAX1 \add_1319/U1_1_13  ( .A(recentdatapoints_len[13]), .B(
        \add_1319/carry[13] ), .YC(\add_1319/carry[14] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[13]) );
  HAX1 \add_1319/U1_1_14  ( .A(recentdatapoints_len[14]), .B(
        \add_1319/carry[14] ), .YC(\add_1319/carry[15] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[14]) );
  HAX1 \add_1319/U1_1_15  ( .A(recentdatapoints_len[15]), .B(
        \add_1319/carry[15] ), .YC(\add_1319/carry[16] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[15]) );
  HAX1 \add_1319/U1_1_16  ( .A(recentdatapoints_len[16]), .B(
        \add_1319/carry[16] ), .YC(\add_1319/carry[17] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[16]) );
  HAX1 \add_1319/U1_1_17  ( .A(recentdatapoints_len[17]), .B(
        \add_1319/carry[17] ), .YC(\add_1319/carry[18] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[17]) );
  HAX1 \add_1319/U1_1_18  ( .A(recentdatapoints_len[18]), .B(
        \add_1319/carry[18] ), .YC(\add_1319/carry[19] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[18]) );
  HAX1 \add_1319/U1_1_19  ( .A(recentdatapoints_len[19]), .B(
        \add_1319/carry[19] ), .YC(\add_1319/carry[20] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[19]) );
  HAX1 \add_1319/U1_1_20  ( .A(recentdatapoints_len[20]), .B(
        \add_1319/carry[20] ), .YC(\add_1319/carry[21] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[20]) );
  HAX1 \add_1319/U1_1_21  ( .A(recentdatapoints_len[21]), .B(
        \add_1319/carry[21] ), .YC(\add_1319/carry[22] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[21]) );
  HAX1 \add_1319/U1_1_22  ( .A(recentdatapoints_len[22]), .B(
        \add_1319/carry[22] ), .YC(\add_1319/carry[23] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[22]) );
  HAX1 \add_1319/U1_1_23  ( .A(recentdatapoints_len[23]), .B(
        \add_1319/carry[23] ), .YC(\add_1319/carry[24] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[23]) );
  HAX1 \add_1319/U1_1_24  ( .A(recentdatapoints_len[24]), .B(
        \add_1319/carry[24] ), .YC(\add_1319/carry[25] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[24]) );
  HAX1 \add_1319/U1_1_25  ( .A(recentdatapoints_len[25]), .B(
        \add_1319/carry[25] ), .YC(\add_1319/carry[26] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[25]) );
  HAX1 \add_1319/U1_1_26  ( .A(recentdatapoints_len[26]), .B(
        \add_1319/carry[26] ), .YC(\add_1319/carry[27] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[26]) );
  HAX1 \add_1319/U1_1_27  ( .A(recentdatapoints_len[27]), .B(
        \add_1319/carry[27] ), .YC(\add_1319/carry[28] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[27]) );
  HAX1 \add_1319/U1_1_28  ( .A(recentdatapoints_len[28]), .B(
        \add_1319/carry[28] ), .YC(\add_1319/carry[29] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[28]) );
  HAX1 \add_1319/U1_1_29  ( .A(recentdatapoints_len[29]), .B(
        \add_1319/carry[29] ), .YC(\add_1319/carry[30] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[29]) );
  HAX1 \add_1319/U1_1_30  ( .A(recentdatapoints_len[30]), .B(
        \add_1319/carry[30] ), .YC(\add_1319/carry[31] ), .YS(
        recentdatapoints_len_load_op_fu_556_p2[30]) );
  FAX1 \sub_1275/U2_1  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[1]), .B(
        n10574), .C(n8648), .YC(\sub_1275/carry[2] ), .YS(i_8_fu_1148_p2[1])
         );
  FAX1 \sub_1275/U2_2  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[2]), .B(
        n10575), .C(\sub_1275/carry[2] ), .YC(\sub_1275/carry[3] ), .YS(
        i_8_fu_1148_p2[2]) );
  FAX1 \sub_1275/U2_3  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[3]), .B(
        n10576), .C(\sub_1275/carry[3] ), .YC(\sub_1275/carry[4] ), .YS(
        i_8_fu_1148_p2[3]) );
  FAX1 \sub_1275/U2_4  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[4]), .B(
        n10577), .C(\sub_1275/carry[4] ), .YC(\sub_1275/carry[5] ), .YS(
        i_8_fu_1148_p2[4]) );
  FAX1 \sub_1275/U2_31  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[31]), 
        .B(n10604), .C(\sub_1275/carry[31] ), .YC(), .YS(i_8_fu_1148_p2[31])
         );
  FAX1 \sub_1269/U2_1  ( .A(CircularBuffer_head_i_read_ass_reg_1624[1]), .B(
        n10140), .C(n8647), .YC(\sub_1269/carry[2] ), .YS(i_5_fu_854_p2[1]) );
  FAX1 \sub_1269/U2_2  ( .A(CircularBuffer_head_i_read_ass_reg_1624[2]), .B(
        n10141), .C(\sub_1269/carry[2] ), .YC(\sub_1269/carry[3] ), .YS(
        i_5_fu_854_p2[2]) );
  FAX1 \sub_1269/U2_3  ( .A(CircularBuffer_head_i_read_ass_reg_1624[3]), .B(
        n10142), .C(\sub_1269/carry[3] ), .YC(\sub_1269/carry[4] ), .YS(
        i_5_fu_854_p2[3]) );
  FAX1 \sub_1269/U2_4  ( .A(CircularBuffer_head_i_read_ass_reg_1624[4]), .B(
        n10143), .C(\sub_1269/carry[4] ), .YC(\sub_1269/carry[5] ), .YS(
        i_5_fu_854_p2[4]) );
  FAX1 \sub_1269/U2_31  ( .A(CircularBuffer_head_i_read_ass_reg_1624[31]), .B(
        n10170), .C(\sub_1269/carry[31] ), .YC(), .YS(i_5_fu_854_p2[31]) );
  FAX1 \sub_1263/U2_1  ( .A(CircularBuffer_head_i_read_ass_reg_1624[1]), .B(
        n10079), .C(n8649), .YC(\sub_1263/carry[2] ), .YS(i_2_fu_823_p2[1]) );
  FAX1 \sub_1263/U2_2  ( .A(CircularBuffer_head_i_read_ass_reg_1624[2]), .B(
        n10080), .C(\sub_1263/carry[2] ), .YC(\sub_1263/carry[3] ), .YS(
        i_2_fu_823_p2[2]) );
  FAX1 \sub_1263/U2_3  ( .A(CircularBuffer_head_i_read_ass_reg_1624[3]), .B(
        n10081), .C(\sub_1263/carry[3] ), .YC(\sub_1263/carry[4] ), .YS(
        i_2_fu_823_p2[3]) );
  FAX1 \sub_1263/U2_4  ( .A(CircularBuffer_head_i_read_ass_reg_1624[4]), .B(
        n10082), .C(\sub_1263/carry[4] ), .YC(\sub_1263/carry[5] ), .YS(
        i_2_fu_823_p2[4]) );
  FAX1 \sub_1263/U2_31  ( .A(CircularBuffer_head_i_read_ass_reg_1624[31]), .B(
        n10109), .C(\sub_1263/carry[31] ), .YC(), .YS(i_2_fu_823_p2[31]) );
  FAX1 \sub_1255/U2_1  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[1]), .B(
        n10635), .C(n8646), .YC(\sub_1255/carry[2] ), .YS(i_11_fu_1179_p2[1])
         );
  FAX1 \sub_1255/U2_2  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[2]), .B(
        n10636), .C(\sub_1255/carry[2] ), .YC(\sub_1255/carry[3] ), .YS(
        i_11_fu_1179_p2[2]) );
  FAX1 \sub_1255/U2_3  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[3]), .B(
        n10637), .C(\sub_1255/carry[3] ), .YC(\sub_1255/carry[4] ), .YS(
        i_11_fu_1179_p2[3]) );
  FAX1 \sub_1255/U2_4  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[4]), .B(
        n10638), .C(\sub_1255/carry[4] ), .YC(\sub_1255/carry[5] ), .YS(
        i_11_fu_1179_p2[4]) );
  FAX1 \sub_1255/U2_31  ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[31]), 
        .B(n10665), .C(\sub_1255/carry[31] ), .YC(), .YS(i_11_fu_1179_p2[31])
         );
  HAX1 \add_1125/U1_1_1  ( .A(recentVBools_len[1]), .B(recentVBools_len[0]), 
        .YC(\add_1125/carry[2] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[1]) );
  HAX1 \add_1125/U1_1_2  ( .A(recentVBools_len[2]), .B(\add_1125/carry[2] ), 
        .YC(\add_1125/carry[3] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[2]) );
  HAX1 \add_1125/U1_1_3  ( .A(recentVBools_len[3]), .B(\add_1125/carry[3] ), 
        .YC(\add_1125/carry[4] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[3]) );
  HAX1 \add_1125/U1_1_4  ( .A(recentVBools_len[4]), .B(\add_1125/carry[4] ), 
        .YC(\add_1125/carry[5] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[4]) );
  HAX1 \add_1125/U1_1_5  ( .A(recentVBools_len[5]), .B(\add_1125/carry[5] ), 
        .YC(\add_1125/carry[6] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[5]) );
  HAX1 \add_1125/U1_1_6  ( .A(recentVBools_len[6]), .B(\add_1125/carry[6] ), 
        .YC(\add_1125/carry[7] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[6]) );
  HAX1 \add_1125/U1_1_7  ( .A(recentVBools_len[7]), .B(\add_1125/carry[7] ), 
        .YC(\add_1125/carry[8] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[7]) );
  HAX1 \add_1125/U1_1_8  ( .A(recentVBools_len[8]), .B(\add_1125/carry[8] ), 
        .YC(\add_1125/carry[9] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[8]) );
  HAX1 \add_1125/U1_1_9  ( .A(recentVBools_len[9]), .B(\add_1125/carry[9] ), 
        .YC(\add_1125/carry[10] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[9]) );
  HAX1 \add_1125/U1_1_10  ( .A(recentVBools_len[10]), .B(\add_1125/carry[10] ), 
        .YC(\add_1125/carry[11] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[10]) );
  HAX1 \add_1125/U1_1_11  ( .A(recentVBools_len[11]), .B(\add_1125/carry[11] ), 
        .YC(\add_1125/carry[12] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[11]) );
  HAX1 \add_1125/U1_1_12  ( .A(recentVBools_len[12]), .B(\add_1125/carry[12] ), 
        .YC(\add_1125/carry[13] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[12]) );
  HAX1 \add_1125/U1_1_13  ( .A(recentVBools_len[13]), .B(\add_1125/carry[13] ), 
        .YC(\add_1125/carry[14] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[13]) );
  HAX1 \add_1125/U1_1_14  ( .A(recentVBools_len[14]), .B(\add_1125/carry[14] ), 
        .YC(\add_1125/carry[15] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[14]) );
  HAX1 \add_1125/U1_1_15  ( .A(recentVBools_len[15]), .B(\add_1125/carry[15] ), 
        .YC(\add_1125/carry[16] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[15]) );
  HAX1 \add_1125/U1_1_16  ( .A(recentVBools_len[16]), .B(\add_1125/carry[16] ), 
        .YC(\add_1125/carry[17] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[16]) );
  HAX1 \add_1125/U1_1_17  ( .A(recentVBools_len[17]), .B(\add_1125/carry[17] ), 
        .YC(\add_1125/carry[18] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[17]) );
  HAX1 \add_1125/U1_1_18  ( .A(recentVBools_len[18]), .B(\add_1125/carry[18] ), 
        .YC(\add_1125/carry[19] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[18]) );
  HAX1 \add_1125/U1_1_19  ( .A(recentVBools_len[19]), .B(\add_1125/carry[19] ), 
        .YC(\add_1125/carry[20] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[19]) );
  HAX1 \add_1125/U1_1_20  ( .A(recentVBools_len[20]), .B(\add_1125/carry[20] ), 
        .YC(\add_1125/carry[21] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[20]) );
  HAX1 \add_1125/U1_1_21  ( .A(recentVBools_len[21]), .B(\add_1125/carry[21] ), 
        .YC(\add_1125/carry[22] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[21]) );
  HAX1 \add_1125/U1_1_22  ( .A(recentVBools_len[22]), .B(\add_1125/carry[22] ), 
        .YC(\add_1125/carry[23] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[22]) );
  HAX1 \add_1125/U1_1_23  ( .A(recentVBools_len[23]), .B(\add_1125/carry[23] ), 
        .YC(\add_1125/carry[24] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[23]) );
  HAX1 \add_1125/U1_1_24  ( .A(recentVBools_len[24]), .B(\add_1125/carry[24] ), 
        .YC(\add_1125/carry[25] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[24]) );
  HAX1 \add_1125/U1_1_25  ( .A(recentVBools_len[25]), .B(\add_1125/carry[25] ), 
        .YC(\add_1125/carry[26] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[25]) );
  HAX1 \add_1125/U1_1_26  ( .A(recentVBools_len[26]), .B(\add_1125/carry[26] ), 
        .YC(\add_1125/carry[27] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[26]) );
  HAX1 \add_1125/U1_1_27  ( .A(recentVBools_len[27]), .B(\add_1125/carry[27] ), 
        .YC(\add_1125/carry[28] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[27]) );
  HAX1 \add_1125/U1_1_28  ( .A(recentVBools_len[28]), .B(\add_1125/carry[28] ), 
        .YC(\add_1125/carry[29] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[28]) );
  HAX1 \add_1125/U1_1_29  ( .A(recentVBools_len[29]), .B(\add_1125/carry[29] ), 
        .YC(\add_1125/carry[30] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[29]) );
  HAX1 \add_1125/U1_1_30  ( .A(recentVBools_len[30]), .B(\add_1125/carry[30] ), 
        .YC(\add_1125/carry[31] ), .YS(
        CircularBuffer_len_read_assign_fu_772_p2[30]) );
  HAX1 \add_1121/U1_1_1  ( .A(recentABools_len[1]), .B(recentABools_len[0]), 
        .YC(\add_1121/carry[2] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[1]) );
  HAX1 \add_1121/U1_1_2  ( .A(recentABools_len[2]), .B(\add_1121/carry[2] ), 
        .YC(\add_1121/carry[3] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[2]) );
  HAX1 \add_1121/U1_1_3  ( .A(recentABools_len[3]), .B(\add_1121/carry[3] ), 
        .YC(\add_1121/carry[4] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[3]) );
  HAX1 \add_1121/U1_1_4  ( .A(recentABools_len[4]), .B(\add_1121/carry[4] ), 
        .YC(\add_1121/carry[5] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[4]) );
  HAX1 \add_1121/U1_1_5  ( .A(recentABools_len[5]), .B(\add_1121/carry[5] ), 
        .YC(\add_1121/carry[6] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[5]) );
  HAX1 \add_1121/U1_1_6  ( .A(recentABools_len[6]), .B(\add_1121/carry[6] ), 
        .YC(\add_1121/carry[7] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[6]) );
  HAX1 \add_1121/U1_1_7  ( .A(recentABools_len[7]), .B(\add_1121/carry[7] ), 
        .YC(\add_1121/carry[8] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[7]) );
  HAX1 \add_1121/U1_1_8  ( .A(recentABools_len[8]), .B(\add_1121/carry[8] ), 
        .YC(\add_1121/carry[9] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[8]) );
  HAX1 \add_1121/U1_1_9  ( .A(recentABools_len[9]), .B(\add_1121/carry[9] ), 
        .YC(\add_1121/carry[10] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[9]) );
  HAX1 \add_1121/U1_1_10  ( .A(recentABools_len[10]), .B(\add_1121/carry[10] ), 
        .YC(\add_1121/carry[11] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[10]) );
  HAX1 \add_1121/U1_1_11  ( .A(recentABools_len[11]), .B(\add_1121/carry[11] ), 
        .YC(\add_1121/carry[12] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[11]) );
  HAX1 \add_1121/U1_1_12  ( .A(recentABools_len[12]), .B(\add_1121/carry[12] ), 
        .YC(\add_1121/carry[13] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[12]) );
  HAX1 \add_1121/U1_1_13  ( .A(recentABools_len[13]), .B(\add_1121/carry[13] ), 
        .YC(\add_1121/carry[14] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[13]) );
  HAX1 \add_1121/U1_1_14  ( .A(recentABools_len[14]), .B(\add_1121/carry[14] ), 
        .YC(\add_1121/carry[15] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[14]) );
  HAX1 \add_1121/U1_1_15  ( .A(recentABools_len[15]), .B(\add_1121/carry[15] ), 
        .YC(\add_1121/carry[16] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[15]) );
  HAX1 \add_1121/U1_1_16  ( .A(recentABools_len[16]), .B(\add_1121/carry[16] ), 
        .YC(\add_1121/carry[17] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[16]) );
  HAX1 \add_1121/U1_1_17  ( .A(recentABools_len[17]), .B(\add_1121/carry[17] ), 
        .YC(\add_1121/carry[18] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[17]) );
  HAX1 \add_1121/U1_1_18  ( .A(recentABools_len[18]), .B(\add_1121/carry[18] ), 
        .YC(\add_1121/carry[19] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[18]) );
  HAX1 \add_1121/U1_1_19  ( .A(recentABools_len[19]), .B(\add_1121/carry[19] ), 
        .YC(\add_1121/carry[20] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[19]) );
  HAX1 \add_1121/U1_1_20  ( .A(recentABools_len[20]), .B(\add_1121/carry[20] ), 
        .YC(\add_1121/carry[21] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[20]) );
  HAX1 \add_1121/U1_1_21  ( .A(recentABools_len[21]), .B(\add_1121/carry[21] ), 
        .YC(\add_1121/carry[22] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[21]) );
  HAX1 \add_1121/U1_1_22  ( .A(recentABools_len[22]), .B(\add_1121/carry[22] ), 
        .YC(\add_1121/carry[23] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[22]) );
  HAX1 \add_1121/U1_1_23  ( .A(recentABools_len[23]), .B(\add_1121/carry[23] ), 
        .YC(\add_1121/carry[24] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[23]) );
  HAX1 \add_1121/U1_1_24  ( .A(recentABools_len[24]), .B(\add_1121/carry[24] ), 
        .YC(\add_1121/carry[25] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[24]) );
  HAX1 \add_1121/U1_1_25  ( .A(recentABools_len[25]), .B(\add_1121/carry[25] ), 
        .YC(\add_1121/carry[26] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[25]) );
  HAX1 \add_1121/U1_1_26  ( .A(recentABools_len[26]), .B(\add_1121/carry[26] ), 
        .YC(\add_1121/carry[27] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[26]) );
  HAX1 \add_1121/U1_1_27  ( .A(recentABools_len[27]), .B(\add_1121/carry[27] ), 
        .YC(\add_1121/carry[28] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[27]) );
  HAX1 \add_1121/U1_1_28  ( .A(recentABools_len[28]), .B(\add_1121/carry[28] ), 
        .YC(\add_1121/carry[29] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[28]) );
  HAX1 \add_1121/U1_1_29  ( .A(recentABools_len[29]), .B(\add_1121/carry[29] ), 
        .YC(\add_1121/carry[30] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[29]) );
  HAX1 \add_1121/U1_1_30  ( .A(recentABools_len[30]), .B(\add_1121/carry[30] ), 
        .YC(\add_1121/carry[31] ), .YS(
        CircularBuffer_len_read_assign_2_fu_1085_p2[30]) );
  AND2X1 U4730 ( .A(n8555), .B(n6349), .Y(n8560) );
  AND2X1 U4731 ( .A(n8549), .B(n7858), .Y(n8552) );
  AND2X1 U4732 ( .A(n8569), .B(n7097), .Y(n8574) );
  AND2X1 U4733 ( .A(n8563), .B(n8387), .Y(n8566) );
  AND2X1 U4734 ( .A(n8554), .B(n6458), .Y(n8558) );
  AND2X1 U4735 ( .A(n8553), .B(n6571), .Y(n8557) );
  AND2X1 U4736 ( .A(n8548), .B(n7640), .Y(n8550) );
  AND2X1 U4737 ( .A(n8557), .B(n6164), .Y(n8559) );
  AND2X1 U4738 ( .A(n8559), .B(n6811), .Y(n8551) );
  AND2X1 U4739 ( .A(n8560), .B(n6686), .Y(n8549) );
  AND2X1 U4740 ( .A(n8552), .B(n7098), .Y(n8556) );
  AND2X1 U4741 ( .A(n8568), .B(n7261), .Y(n8572) );
  AND2X1 U4742 ( .A(n8567), .B(n7435), .Y(n8571) );
  AND2X1 U4743 ( .A(n8562), .B(n8101), .Y(n8564) );
  AND2X1 U4744 ( .A(n8571), .B(n7096), .Y(n8573) );
  AND2X1 U4745 ( .A(n8573), .B(n7436), .Y(n8565) );
  AND2X1 U4746 ( .A(n8574), .B(n7262), .Y(n8563) );
  OR2X1 U4747 ( .A(n6800), .B(n6799), .Y(n2050) );
  AND2X1 U4748 ( .A(n8566), .B(n7639), .Y(n8570) );
  AND2X1 U4749 ( .A(n7833), .B(sum_1_phi_fu_379_p4[30]), .Y(n11778) );
  AND2X1 U4750 ( .A(n6019), .B(n4692), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n362 )
         );
  AND2X1 U4751 ( .A(n6951), .B(n6952), .Y(n11081) );
  AND2X1 U4752 ( .A(n8107), .B(n6093), .Y(n8554) );
  AND2X1 U4753 ( .A(n8558), .B(n6946), .Y(n8548) );
  AND2X1 U4754 ( .A(n8550), .B(n7437), .Y(n8553) );
  AND2X1 U4755 ( .A(n8551), .B(n7263), .Y(n8555) );
  AND2X1 U4756 ( .A(n8556), .B(n6252), .Y(n8561) );
  AND2X1 U4757 ( .A(n7832), .B(sum_phi_fu_311_p4[30]), .Y(n11520) );
  AND2X1 U4758 ( .A(n8390), .B(n6944), .Y(n8568) );
  AND2X1 U4759 ( .A(n8572), .B(n7638), .Y(n8562) );
  AND2X1 U4760 ( .A(n8564), .B(n7857), .Y(n8567) );
  AND2X1 U4761 ( .A(n8565), .B(n7856), .Y(n8569) );
  AND2X1 U4762 ( .A(n8570), .B(n6945), .Y(n8575) );
  AND2X1 U4763 ( .A(n6951), .B(n6952), .Y(n11063) );
  AND2X1 U4764 ( .A(n7586), .B(n11617), .Y(n11619) );
  AND2X1 U4765 ( .A(n8561), .B(n8408), .Y(n8636) );
  AND2X1 U4766 ( .A(n7584), .B(n12250), .Y(n12252) );
  AND2X1 U4767 ( .A(n8575), .B(n8115), .Y(n8637) );
  AND2X1 U4768 ( .A(n8888), .B(n6018), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n352 )
         );
  AND2X1 U4769 ( .A(n6019), .B(n9823), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n354 )
         );
  OR2X1 U4770 ( .A(n8857), .B(n8268), .Y(\Decision_AXILiteS_s_axi_U/n332 ) );
  AND2X1 U4771 ( .A(n4696), .B(n9481), .Y(n11573) );
  AND2X1 U4772 ( .A(n4697), .B(n4774), .Y(n11622) );
  AND2X1 U4773 ( .A(n4698), .B(n9498), .Y(n12206) );
  AND2X1 U4774 ( .A(n4699), .B(n4775), .Y(n12255) );
  AND2X1 U4775 ( .A(n7588), .B(n10449), .Y(n11916) );
  OR2X1 U4776 ( .A(n6679), .B(recentABools_data_address0[3]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n31 ) );
  OR2X1 U4777 ( .A(n7404), .B(recentVBools_data_address0[3]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n25 ) );
  OR2X1 U4778 ( .A(n6678), .B(recentVBools_data_address0[3]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n30 ) );
  OR2X1 U4779 ( .A(n5226), .B(n8100), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n13 ) );
  OR2X1 U4780 ( .A(n5225), .B(n8100), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n8 ) );
  AND2X1 U4781 ( .A(n8889), .B(n6012), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 )
         );
  AND2X1 U4782 ( .A(n6012), .B(n9822), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 )
         );
  OR2X1 U4783 ( .A(n7847), .B(\Decision_AXILiteS_s_axi_U/waddr[2] ), .Y(
        \Decision_AXILiteS_s_axi_U/n576 ) );
  OR2X1 U4784 ( .A(n8394), .B(n8395), .Y(\toReturn_1_fu_1395_p3[7] ) );
  AND2X1 U4785 ( .A(n11194), .B(n6166), .Y(n11196) );
  AND2X1 U4786 ( .A(n11224), .B(n6165), .Y(n11226) );
  OR2X1 U4787 ( .A(n5259), .B(n5292), .Y(n1928) );
  OR2X1 U4788 ( .A(n8380), .B(n8381), .Y(n2018) );
  OR2X1 U4789 ( .A(n5258), .B(n5291), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n342 )
         );
  OR2X1 U4790 ( .A(n5257), .B(n5290), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n343 )
         );
  OR2X1 U4791 ( .A(n5256), .B(n5289), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n321 )
         );
  OR2X1 U4792 ( .A(n5255), .B(n5288), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n322 )
         );
  OR2X1 U4793 ( .A(n5254), .B(n5287), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n300 )
         );
  OR2X1 U4794 ( .A(n5253), .B(n5286), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n301 )
         );
  OR2X1 U4795 ( .A(n5252), .B(n5285), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n279 )
         );
  OR2X1 U4796 ( .A(n5251), .B(n5284), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n280 )
         );
  OR2X1 U4797 ( .A(n5250), .B(n5283), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n258 )
         );
  OR2X1 U4798 ( .A(n5249), .B(n5282), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n259 )
         );
  OR2X1 U4799 ( .A(n5248), .B(n5281), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n237 )
         );
  OR2X1 U4800 ( .A(n5247), .B(n5280), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n238 )
         );
  OR2X1 U4801 ( .A(n5246), .B(n5279), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n216 )
         );
  OR2X1 U4802 ( .A(n5245), .B(n5278), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n217 )
         );
  OR2X1 U4803 ( .A(n5244), .B(n5277), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n195 )
         );
  OR2X1 U4804 ( .A(n5243), .B(n5276), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n196 )
         );
  OR2X1 U4805 ( .A(n5242), .B(n5275), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n174 )
         );
  OR2X1 U4806 ( .A(n5241), .B(n5274), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n175 )
         );
  OR2X1 U4807 ( .A(n5240), .B(n5273), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n153 )
         );
  OR2X1 U4808 ( .A(n5239), .B(n5272), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n154 )
         );
  OR2X1 U4809 ( .A(n5238), .B(n5271), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n132 )
         );
  OR2X1 U4810 ( .A(n5237), .B(n5270), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n133 )
         );
  OR2X1 U4811 ( .A(n5236), .B(n5269), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n111 )
         );
  OR2X1 U4812 ( .A(n5235), .B(n5268), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n112 )
         );
  OR2X1 U4813 ( .A(n5234), .B(n5267), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n90 ) );
  OR2X1 U4814 ( .A(n5233), .B(n5266), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n91 ) );
  OR2X1 U4815 ( .A(n5232), .B(n5265), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n69 ) );
  OR2X1 U4816 ( .A(n5231), .B(n5264), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n70 ) );
  OR2X1 U4817 ( .A(n5230), .B(n5263), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n48 ) );
  OR2X1 U4818 ( .A(n5229), .B(n5262), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n49 ) );
  OR2X1 U4819 ( .A(n5228), .B(n5261), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n5 ) );
  OR2X1 U4820 ( .A(n5227), .B(n5260), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n6 ) );
  AND2X1 U4821 ( .A(ap_rst_n), .B(n4794), .Y(\Decision_AXILiteS_s_axi_U/n612 )
         );
  AND2X1 U4822 ( .A(ap_rst_n), .B(n8106), .Y(\Decision_AXILiteS_s_axi_U/n607 )
         );
  AND2X1 U4823 ( .A(ap_rst_n), .B(n8412), .Y(\Decision_AXILiteS_s_axi_U/n462 )
         );
  AND2X1 U4824 ( .A(n8411), .B(\Decision_AXILiteS_s_axi_U/n565 ), .Y(
        \Decision_AXILiteS_s_axi_U/n460 ) );
  AND2X1 U4825 ( .A(n4708), .B(n4784), .Y(\Decision_AXILiteS_s_axi_U/n252 ) );
  AND2X1 U4826 ( .A(n4709), .B(n4785), .Y(\Decision_AXILiteS_s_axi_U/n262 ) );
  AND2X1 U4827 ( .A(n4710), .B(n4786), .Y(\Decision_AXILiteS_s_axi_U/n269 ) );
  AND2X1 U4828 ( .A(n4711), .B(n4787), .Y(\Decision_AXILiteS_s_axi_U/n276 ) );
  AND2X1 U4829 ( .A(n4712), .B(n4788), .Y(\Decision_AXILiteS_s_axi_U/n282 ) );
  AND2X1 U4830 ( .A(n4713), .B(n4789), .Y(\Decision_AXILiteS_s_axi_U/n291 ) );
  AND2X1 U4831 ( .A(ap_rst_n), .B(n7083), .Y(n8427) );
  OR2X1 U4832 ( .A(n8386), .B(n2238), .Y(n11197) );
  OR2X1 U4833 ( .A(n8385), .B(n2734), .Y(n11227) );
  AND2X1 U4834 ( .A(ap_rst_n), .B(n4793), .Y(\Decision_AXILiteS_s_axi_U/n572 )
         );
  AND2X1 U4835 ( .A(ap_rst_n), .B(n4792), .Y(\Decision_AXILiteS_s_axi_U/n567 )
         );
  AND2X1 U4836 ( .A(n4700), .B(n4776), .Y(\Decision_AXILiteS_s_axi_U/n207 ) );
  AND2X1 U4837 ( .A(n4701), .B(n4777), .Y(\Decision_AXILiteS_s_axi_U/n214 ) );
  AND2X1 U4838 ( .A(n4702), .B(n4778), .Y(\Decision_AXILiteS_s_axi_U/n219 ) );
  AND2X1 U4839 ( .A(n4703), .B(n4779), .Y(\Decision_AXILiteS_s_axi_U/n224 ) );
  AND2X1 U4840 ( .A(n4704), .B(n4780), .Y(\Decision_AXILiteS_s_axi_U/n229 ) );
  AND2X1 U4841 ( .A(n4705), .B(n4781), .Y(\Decision_AXILiteS_s_axi_U/n234 ) );
  AND2X1 U4842 ( .A(n4706), .B(n4782), .Y(\Decision_AXILiteS_s_axi_U/n239 ) );
  AND2X1 U4843 ( .A(n4707), .B(n4783), .Y(\Decision_AXILiteS_s_axi_U/n244 ) );
  AND2X1 U4844 ( .A(n8306), .B(n7982), .Y(n3650) );
  AND2X1 U4845 ( .A(n8062), .B(n7764), .Y(n3653) );
  AND2X1 U4846 ( .A(n7840), .B(n7566), .Y(n3656) );
  AND2X1 U4847 ( .A(n7628), .B(n7385), .Y(n3659) );
  AND2X1 U4848 ( .A(n8222), .B(n8223), .Y(n3783) );
  AND2X1 U4849 ( .A(n8305), .B(n7980), .Y(n3854) );
  AND2X1 U4850 ( .A(n8061), .B(n7762), .Y(n3857) );
  AND2X1 U4851 ( .A(n7627), .B(n7383), .Y(n3858) );
  AND2X1 U4852 ( .A(n7839), .B(n7564), .Y(n3861) );
  AND2X1 U4853 ( .A(n7997), .B(n7996), .Y(n4539) );
  AND2X1 U4854 ( .A(n8235), .B(n8234), .Y(n4540) );
  AND2X1 U4855 ( .A(n7776), .B(n7775), .Y(n4541) );
  AND2X1 U4856 ( .A(n7582), .B(n7581), .Y(n4542) );
  AND2X1 U4857 ( .A(n7397), .B(n7396), .Y(n4543) );
  AND2X1 U4858 ( .A(n7232), .B(n7231), .Y(n4544) );
  AND2X1 U4859 ( .A(n7076), .B(n7075), .Y(n4545) );
  AND2X1 U4860 ( .A(n6933), .B(n6932), .Y(n4546) );
  AND2X1 U4861 ( .A(n6798), .B(n6797), .Y(n4547) );
  AND2X1 U4862 ( .A(n6677), .B(n6676), .Y(n4548) );
  AND2X1 U4863 ( .A(n6568), .B(n6567), .Y(n4549) );
  AND2X1 U4864 ( .A(n6455), .B(n6454), .Y(n4550) );
  AND2X1 U4865 ( .A(n7994), .B(n7993), .Y(n4551) );
  AND2X1 U4866 ( .A(n6346), .B(n6345), .Y(n4552) );
  AND2X1 U4867 ( .A(n6251), .B(n6250), .Y(n4553) );
  AND2X1 U4868 ( .A(n6163), .B(n6162), .Y(n4554) );
  AND2X1 U4869 ( .A(n7579), .B(n7578), .Y(n4555) );
  AND2X1 U4870 ( .A(n8232), .B(n8231), .Y(n4556) );
  AND2X1 U4871 ( .A(n7773), .B(n7772), .Y(n4557) );
  AND2X1 U4872 ( .A(n7394), .B(n7393), .Y(n4558) );
  AND2X1 U4873 ( .A(n7229), .B(n7228), .Y(n4559) );
  AND2X1 U4874 ( .A(n7073), .B(n7072), .Y(n4560) );
  AND2X1 U4875 ( .A(n6930), .B(n6929), .Y(n4561) );
  AND2X1 U4876 ( .A(n6795), .B(n6794), .Y(n4562) );
  AND2X1 U4877 ( .A(n6674), .B(n6673), .Y(n4563) );
  AND2X1 U4878 ( .A(n7991), .B(n7990), .Y(n4564) );
  AND2X1 U4879 ( .A(n6565), .B(n6564), .Y(n4565) );
  AND2X1 U4880 ( .A(n6452), .B(n6451), .Y(n4566) );
  AND2X1 U4881 ( .A(n6343), .B(n6342), .Y(n4567) );
  AND2X1 U4882 ( .A(n6248), .B(n6247), .Y(n4568) );
  AND2X1 U4883 ( .A(n8229), .B(n8228), .Y(n4569) );
  AND2X1 U4884 ( .A(n7770), .B(n7769), .Y(n4570) );
  AND2X1 U4885 ( .A(n7576), .B(n7575), .Y(n4603) );
  AND2X1 U4886 ( .A(n7391), .B(n7390), .Y(n4604) );
  AND2X1 U4887 ( .A(n7226), .B(n7225), .Y(n4605) );
  AND2X1 U4888 ( .A(n7070), .B(n7069), .Y(n4606) );
  AND2X1 U4889 ( .A(n6927), .B(n6926), .Y(n4607) );
  AND2X1 U4890 ( .A(n6792), .B(n6791), .Y(n4608) );
  AND2X1 U4891 ( .A(n7988), .B(n7987), .Y(n4609) );
  AND2X1 U4892 ( .A(n6671), .B(n6670), .Y(n4610) );
  AND2X1 U4893 ( .A(n6562), .B(n6561), .Y(n4611) );
  AND2X1 U4894 ( .A(n6449), .B(n6448), .Y(n4612) );
  AND2X1 U4895 ( .A(n6340), .B(n6339), .Y(n4613) );
  AND2X1 U4896 ( .A(n6245), .B(n6244), .Y(n4614) );
  AND2X1 U4897 ( .A(n6160), .B(n6159), .Y(n4615) );
  AND2X1 U4898 ( .A(n8226), .B(n8225), .Y(n4616) );
  AND2X1 U4899 ( .A(n7767), .B(n7766), .Y(n4617) );
  AND2X1 U4900 ( .A(n7573), .B(n7572), .Y(n4618) );
  AND2X1 U4901 ( .A(n7388), .B(n7387), .Y(n4619) );
  AND2X1 U4902 ( .A(n7223), .B(n7222), .Y(n4620) );
  AND2X1 U4903 ( .A(n7067), .B(n7066), .Y(n4621) );
  AND2X1 U4904 ( .A(n7985), .B(n7984), .Y(n4622) );
  AND2X1 U4905 ( .A(n6924), .B(n6923), .Y(n4623) );
  AND2X1 U4906 ( .A(n6789), .B(n6788), .Y(n4624) );
  AND2X1 U4907 ( .A(n6157), .B(n6156), .Y(n4625) );
  AND2X1 U4908 ( .A(n6668), .B(n6667), .Y(n4626) );
  AND2X1 U4909 ( .A(n6559), .B(n6558), .Y(n4627) );
  AND2X1 U4910 ( .A(n6446), .B(n6445), .Y(n4628) );
  AND2X1 U4911 ( .A(n6337), .B(n6336), .Y(n4629) );
  AND2X1 U4912 ( .A(n6242), .B(n6241), .Y(n4630) );
  AND2X1 U4913 ( .A(n6088), .B(n6087), .Y(n4631) );
  AND2X1 U4914 ( .A(n8219), .B(n8220), .Y(n4054) );
  AND2X1 U4915 ( .A(n4714), .B(n4790), .Y(recentABools_data_address0[4]) );
  AND2X1 U4916 ( .A(n4715), .B(n4791), .Y(recentVBools_data_address0[4]) );
  AND2X1 U4917 ( .A(ap_CS_fsm[1]), .B(n8294), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ) );
  AND2X1 U4918 ( .A(n7649), .B(n7650), .Y(recentABools_data_address0[2]) );
  AND2X1 U4919 ( .A(n8414), .B(n8415), .Y(recentVBools_data_address0[2]) );
  AND2X1 U4920 ( .A(n6802), .B(n6801), .Y(n8644) );
  AND2X1 U4921 ( .A(n6804), .B(n6803), .Y(n8645) );
  AND2X1 U4922 ( .A(n2533), .B(n8378), .Y(n2535) );
  AND2X1 U4923 ( .A(n7254), .B(n7253), .Y(recentABools_data_address0[0]) );
  AND2X1 U4924 ( .A(n7430), .B(n7429), .Y(recentVBools_data_address0[0]) );
  OR2X1 U4925 ( .A(n8978), .B(n8379), .Y(n8428) );
  XNOR2X1 U4926 ( .A(CircularBuffer_int_30_sum_i_fu_758_p3[31]), .B(n8855), 
        .Y(n4688) );
  XNOR2X1 U4927 ( .A(CircularBuffer_int_30_sum_i1_fu_1071_p3[31]), .B(n8856), 
        .Y(n4689) );
  OR2X1 U4928 ( .A(n6090), .B(n6089), .Y(n3151) );
  OR2X1 U4929 ( .A(n6092), .B(n6091), .Y(n3149) );
  AND2X1 U4930 ( .A(n8927), .B(n8293), .Y(n2701) );
  AND2X1 U4931 ( .A(n8934), .B(n8292), .Y(n2241) );
  AND2X1 U4932 ( .A(n8109), .B(n8110), .Y(recentVBools_data_address0[3]) );
  AND2X1 U4933 ( .A(n8403), .B(n8404), .Y(recentABools_data_address0[3]) );
  AND2X1 U4934 ( .A(ap_rst_n), .B(n7842), .Y(n8429) );
  OR2X1 U4935 ( .A(n5713), .B(n5714), .Y(n5712) );
  OR2X1 U4936 ( .A(n5854), .B(\Decision_AXILiteS_s_axi_U/n302 ), .Y(n5714) );
  OR2X1 U4937 ( .A(n5716), .B(n5717), .Y(n5715) );
  OR2X1 U4938 ( .A(n5857), .B(\Decision_AXILiteS_s_axi_U/n317 ), .Y(n5717) );
  OR2X1 U4939 ( .A(n5956), .B(n5944), .Y(n5942) );
  INVX1 U4940 ( .A(n5942), .Y(n4690) );
  OR2X1 U4941 ( .A(n5943), .B(n11563), .Y(n5944) );
  OR2X1 U4942 ( .A(n5959), .B(n5947), .Y(n5945) );
  INVX1 U4943 ( .A(n5945), .Y(n4691) );
  OR2X1 U4944 ( .A(n5946), .B(n12196), .Y(n5947) );
  OR2X1 U4945 ( .A(n11559), .B(n5958), .Y(n5956) );
  OR2X1 U4946 ( .A(n5957), .B(n11558), .Y(n5958) );
  OR2X1 U4947 ( .A(n12192), .B(n5961), .Y(n5959) );
  OR2X1 U4948 ( .A(n5960), .B(n12191), .Y(n5961) );
  OR2X1 U4949 ( .A(n5973), .B(n5974), .Y(n5971) );
  OR2X1 U4950 ( .A(n5972), .B(n346), .Y(n5974) );
  OR2X1 U4951 ( .A(n6014), .B(n6015), .Y(n6012) );
  INVX1 U4952 ( .A(n6012), .Y(n4692) );
  OR2X1 U4953 ( .A(n6013), .B(n356), .Y(n6015) );
  OR2X1 U4954 ( .A(n6021), .B(n6022), .Y(n6019) );
  INVX1 U4955 ( .A(n6019), .Y(n4693) );
  OR2X1 U4956 ( .A(n6020), .B(n353), .Y(n6022) );
  OR2X1 U4957 ( .A(recentABools_data_address0[4]), .B(n6026), .Y(n6024) );
  INVX1 U4958 ( .A(n6024), .Y(n4694) );
  OR2X1 U4959 ( .A(n6025), .B(recentABools_data_address0[3]), .Y(n6026) );
  OR2X1 U4960 ( .A(recentVBools_data_address0[4]), .B(n6029), .Y(n6027) );
  INVX1 U4961 ( .A(n6027), .Y(n4695) );
  OR2X1 U4962 ( .A(n6028), .B(recentVBools_data_address0[3]), .Y(n6029) );
  AND2X1 U4963 ( .A(n8547), .B(CircularBuffer_int_30_sum_i_fu_758_p3[30]), .Y(
        n8855) );
  AND2X1 U4964 ( .A(n8546), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[30]), 
        .Y(n8856) );
  AND2X1 U4965 ( .A(a_thresh[29]), .B(n9490), .Y(n11559) );
  AND2X1 U4966 ( .A(a_thresh[28]), .B(n9490), .Y(n11558) );
  AND2X1 U4967 ( .A(a_thresh[25]), .B(n9490), .Y(n11563) );
  AND2X1 U4968 ( .A(v_thresh[29]), .B(n9540), .Y(n12192) );
  AND2X1 U4969 ( .A(v_thresh[28]), .B(n9540), .Y(n12191) );
  AND2X1 U4970 ( .A(v_thresh[25]), .B(n9540), .Y(n12196) );
  AND2X1 U4971 ( .A(v_flip[1]), .B(n9314), .Y(\Decision_AXILiteS_s_axi_U/n302 ) );
  AND2X1 U4972 ( .A(v_flip[0]), .B(n9314), .Y(\Decision_AXILiteS_s_axi_U/n317 ) );
  OR2X1 U4973 ( .A(n8968), .B(\reset_params_V[0] ), .Y(n2872) );
  AND2X1 U4974 ( .A(i_fu_607_p2[2]), .B(n349), .Y(n356) );
  AND2X1 U4975 ( .A(i_fu_607_p2[3]), .B(n349), .Y(n353) );
  AND2X1 U4976 ( .A(i_fu_607_p2[4]), .B(n349), .Y(n346) );
  BUFX2 U4977 ( .A(n11568), .Y(n4696) );
  BUFX2 U4978 ( .A(n11614), .Y(n4697) );
  BUFX2 U4979 ( .A(n12201), .Y(n4698) );
  BUFX2 U4980 ( .A(n12247), .Y(n4699) );
  BUFX2 U4981 ( .A(\Decision_AXILiteS_s_axi_U/n208 ), .Y(n4700) );
  BUFX2 U4982 ( .A(\Decision_AXILiteS_s_axi_U/n215 ), .Y(n4701) );
  BUFX2 U4983 ( .A(\Decision_AXILiteS_s_axi_U/n220 ), .Y(n4702) );
  BUFX2 U4984 ( .A(\Decision_AXILiteS_s_axi_U/n225 ), .Y(n4703) );
  BUFX2 U4985 ( .A(\Decision_AXILiteS_s_axi_U/n230 ), .Y(n4704) );
  BUFX2 U4986 ( .A(\Decision_AXILiteS_s_axi_U/n235 ), .Y(n4705) );
  BUFX2 U4987 ( .A(\Decision_AXILiteS_s_axi_U/n240 ), .Y(n4706) );
  BUFX2 U4988 ( .A(\Decision_AXILiteS_s_axi_U/n245 ), .Y(n4707) );
  BUFX2 U4989 ( .A(\Decision_AXILiteS_s_axi_U/n253 ), .Y(n4708) );
  BUFX2 U4990 ( .A(\Decision_AXILiteS_s_axi_U/n263 ), .Y(n4709) );
  BUFX2 U4991 ( .A(\Decision_AXILiteS_s_axi_U/n270 ), .Y(n4710) );
  BUFX2 U4992 ( .A(\Decision_AXILiteS_s_axi_U/n277 ), .Y(n4711) );
  BUFX2 U4993 ( .A(\Decision_AXILiteS_s_axi_U/n283 ), .Y(n4712) );
  BUFX2 U4994 ( .A(\Decision_AXILiteS_s_axi_U/n292 ), .Y(n4713) );
  BUFX2 U4995 ( .A(n383), .Y(n4714) );
  BUFX2 U4996 ( .A(n369), .Y(n4715) );
  BUFX2 U4997 ( .A(n3785), .Y(n4716) );
  BUFX2 U4998 ( .A(n3452), .Y(n4717) );
  BUFX2 U4999 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n893 ), 
        .Y(n4718) );
  BUFX2 U5000 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n894 ), 
        .Y(n4719) );
  BUFX2 U5001 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n895 ), 
        .Y(n4720) );
  BUFX2 U5002 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n896 ), 
        .Y(n4721) );
  BUFX2 U5003 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n897 ), 
        .Y(n4722) );
  BUFX2 U5004 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n898 ), 
        .Y(n4723) );
  BUFX2 U5005 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n899 ), 
        .Y(n4724) );
  BUFX2 U5006 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n900 ), 
        .Y(n4725) );
  BUFX2 U5007 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n901 ), 
        .Y(n4726) );
  BUFX2 U5008 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n902 ), 
        .Y(n4727) );
  BUFX2 U5009 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n903 ), 
        .Y(n4728) );
  BUFX2 U5010 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n904 ), 
        .Y(n4729) );
  BUFX2 U5011 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n905 ), 
        .Y(n4730) );
  BUFX2 U5012 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n906 ), 
        .Y(n4731) );
  BUFX2 U5013 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n907 ), 
        .Y(n4732) );
  BUFX2 U5014 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n908 ), 
        .Y(n4733) );
  BUFX2 U5015 ( .A(\Decision_AXILiteS_s_axi_U/n648 ), .Y(n4734) );
  BUFX2 U5016 ( .A(\Decision_AXILiteS_s_axi_U/n649 ), .Y(n4735) );
  BUFX2 U5017 ( .A(\Decision_AXILiteS_s_axi_U/n650 ), .Y(n4736) );
  BUFX2 U5018 ( .A(\Decision_AXILiteS_s_axi_U/n651 ), .Y(n4737) );
  BUFX2 U5019 ( .A(\Decision_AXILiteS_s_axi_U/n652 ), .Y(n4738) );
  BUFX2 U5020 ( .A(\Decision_AXILiteS_s_axi_U/n653 ), .Y(n4739) );
  BUFX2 U5021 ( .A(\Decision_AXILiteS_s_axi_U/n654 ), .Y(n4740) );
  BUFX2 U5022 ( .A(\Decision_AXILiteS_s_axi_U/n655 ), .Y(n4741) );
  BUFX2 U5023 ( .A(\Decision_AXILiteS_s_axi_U/n656 ), .Y(n4742) );
  BUFX2 U5024 ( .A(\Decision_AXILiteS_s_axi_U/n657 ), .Y(n4743) );
  BUFX2 U5025 ( .A(\Decision_AXILiteS_s_axi_U/n658 ), .Y(n4744) );
  BUFX2 U5026 ( .A(\Decision_AXILiteS_s_axi_U/n659 ), .Y(n4745) );
  BUFX2 U5027 ( .A(\Decision_AXILiteS_s_axi_U/n660 ), .Y(n4746) );
  BUFX2 U5028 ( .A(\Decision_AXILiteS_s_axi_U/n661 ), .Y(n4747) );
  BUFX2 U5029 ( .A(\Decision_AXILiteS_s_axi_U/n662 ), .Y(n4748) );
  BUFX2 U5030 ( .A(\Decision_AXILiteS_s_axi_U/n663 ), .Y(n4749) );
  BUFX2 U5031 ( .A(\Decision_AXILiteS_s_axi_U/n664 ), .Y(n4750) );
  BUFX2 U5032 ( .A(\Decision_AXILiteS_s_axi_U/n665 ), .Y(n4751) );
  BUFX2 U5033 ( .A(\Decision_AXILiteS_s_axi_U/n666 ), .Y(n4752) );
  BUFX2 U5034 ( .A(\Decision_AXILiteS_s_axi_U/n667 ), .Y(n4753) );
  BUFX2 U5035 ( .A(\Decision_AXILiteS_s_axi_U/n668 ), .Y(n4754) );
  BUFX2 U5036 ( .A(\Decision_AXILiteS_s_axi_U/n669 ), .Y(n4755) );
  BUFX2 U5037 ( .A(\Decision_AXILiteS_s_axi_U/n670 ), .Y(n4756) );
  BUFX2 U5038 ( .A(\Decision_AXILiteS_s_axi_U/n671 ), .Y(n4757) );
  BUFX2 U5039 ( .A(\Decision_AXILiteS_s_axi_U/n856 ), .Y(n4758) );
  BUFX2 U5040 ( .A(N105), .Y(n4759) );
  BUFX2 U5041 ( .A(N110), .Y(n4760) );
  BUFX2 U5042 ( .A(N98), .Y(n4761) );
  AND2X1 U5043 ( .A(n5219), .B(n5199), .Y(\Decision_AXILiteS_s_axi_U/n873 ) );
  INVX1 U5044 ( .A(\Decision_AXILiteS_s_axi_U/n873 ), .Y(n4762) );
  AND2X1 U5045 ( .A(n5216), .B(n5200), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n88 ) );
  INVX1 U5046 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n88 ), 
        .Y(n4763) );
  AND2X1 U5047 ( .A(n5217), .B(n5201), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n86 ) );
  INVX1 U5048 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n86 ), 
        .Y(n4764) );
  AND2X1 U5049 ( .A(n5220), .B(\Decision_AXILiteS_s_axi_U/n250 ), .Y(
        \Decision_AXILiteS_s_axi_U/n672 ) );
  INVX1 U5050 ( .A(\Decision_AXILiteS_s_axi_U/n672 ), .Y(n4765) );
  AND2X1 U5051 ( .A(n5221), .B(\Decision_AXILiteS_s_axi_U/n280 ), .Y(
        \Decision_AXILiteS_s_axi_U/n673 ) );
  INVX1 U5052 ( .A(\Decision_AXILiteS_s_axi_U/n673 ), .Y(n4766) );
  AND2X1 U5053 ( .A(n5222), .B(\Decision_AXILiteS_s_axi_U/n289 ), .Y(
        \Decision_AXILiteS_s_axi_U/n674 ) );
  INVX1 U5054 ( .A(\Decision_AXILiteS_s_axi_U/n674 ), .Y(n4767) );
  AND2X1 U5055 ( .A(n5223), .B(\Decision_AXILiteS_s_axi_U/n298 ), .Y(
        \Decision_AXILiteS_s_axi_U/n675 ) );
  INVX1 U5056 ( .A(\Decision_AXILiteS_s_axi_U/n675 ), .Y(n4768) );
  AND2X1 U5057 ( .A(n5224), .B(\Decision_AXILiteS_s_axi_U/n312 ), .Y(
        \Decision_AXILiteS_s_axi_U/n676 ) );
  INVX1 U5058 ( .A(\Decision_AXILiteS_s_axi_U/n676 ), .Y(n4769) );
  AND2X1 U5059 ( .A(n5218), .B(n7842), .Y(\Decision_AXILiteS_s_axi_U/n863 ) );
  INVX1 U5060 ( .A(\Decision_AXILiteS_s_axi_U/n863 ), .Y(n4770) );
  AND2X1 U5061 ( .A(n5205), .B(n5202), .Y(n4634) );
  INVX1 U5062 ( .A(n4634), .Y(n4771) );
  AND2X1 U5063 ( .A(n5206), .B(n5203), .Y(n4633) );
  INVX1 U5064 ( .A(n4633), .Y(n4772) );
  AND2X1 U5065 ( .A(n5207), .B(n5204), .Y(n4632) );
  INVX1 U5066 ( .A(n4632), .Y(n4773) );
  BUFX2 U5067 ( .A(n11613), .Y(n4774) );
  BUFX2 U5068 ( .A(n12246), .Y(n4775) );
  BUFX2 U5069 ( .A(\Decision_AXILiteS_s_axi_U/n209 ), .Y(n4776) );
  BUFX2 U5070 ( .A(\Decision_AXILiteS_s_axi_U/n216 ), .Y(n4777) );
  BUFX2 U5071 ( .A(\Decision_AXILiteS_s_axi_U/n221 ), .Y(n4778) );
  BUFX2 U5072 ( .A(\Decision_AXILiteS_s_axi_U/n226 ), .Y(n4779) );
  BUFX2 U5073 ( .A(\Decision_AXILiteS_s_axi_U/n231 ), .Y(n4780) );
  BUFX2 U5074 ( .A(\Decision_AXILiteS_s_axi_U/n236 ), .Y(n4781) );
  BUFX2 U5075 ( .A(\Decision_AXILiteS_s_axi_U/n241 ), .Y(n4782) );
  BUFX2 U5076 ( .A(\Decision_AXILiteS_s_axi_U/n246 ), .Y(n4783) );
  BUFX2 U5077 ( .A(\Decision_AXILiteS_s_axi_U/n254 ), .Y(n4784) );
  BUFX2 U5078 ( .A(\Decision_AXILiteS_s_axi_U/n264 ), .Y(n4785) );
  BUFX2 U5079 ( .A(\Decision_AXILiteS_s_axi_U/n271 ), .Y(n4786) );
  BUFX2 U5080 ( .A(\Decision_AXILiteS_s_axi_U/n278 ), .Y(n4787) );
  BUFX2 U5081 ( .A(\Decision_AXILiteS_s_axi_U/n284 ), .Y(n4788) );
  BUFX2 U5082 ( .A(\Decision_AXILiteS_s_axi_U/n293 ), .Y(n4789) );
  BUFX2 U5083 ( .A(n384), .Y(n4790) );
  BUFX2 U5084 ( .A(n370), .Y(n4791) );
  BUFX2 U5085 ( .A(\Decision_AXILiteS_s_axi_U/n569 ), .Y(n4792) );
  BUFX2 U5086 ( .A(\Decision_AXILiteS_s_axi_U/n574 ), .Y(n4793) );
  BUFX2 U5087 ( .A(\Decision_AXILiteS_s_axi_U/n614 ), .Y(n4794) );
  BUFX2 U5088 ( .A(n2863), .Y(n4795) );
  BUFX2 U5089 ( .A(n2861), .Y(n4796) );
  BUFX2 U5090 ( .A(n2763), .Y(n4797) );
  BUFX2 U5091 ( .A(n2761), .Y(n4798) );
  BUFX2 U5092 ( .A(n2755), .Y(n4799) );
  BUFX2 U5093 ( .A(n2753), .Y(n4800) );
  BUFX2 U5094 ( .A(n2751), .Y(n4801) );
  BUFX2 U5095 ( .A(n2739), .Y(n4802) );
  BUFX2 U5096 ( .A(n2737), .Y(n4803) );
  BUFX2 U5097 ( .A(n2402), .Y(n4804) );
  BUFX2 U5098 ( .A(n2400), .Y(n4805) );
  BUFX2 U5099 ( .A(n2278), .Y(n4806) );
  BUFX2 U5100 ( .A(n2276), .Y(n4807) );
  BUFX2 U5101 ( .A(n2270), .Y(n4808) );
  BUFX2 U5102 ( .A(n2268), .Y(n4809) );
  BUFX2 U5103 ( .A(n2266), .Y(n4810) );
  BUFX2 U5104 ( .A(n2262), .Y(n4811) );
  BUFX2 U5105 ( .A(n2260), .Y(n4812) );
  BUFX2 U5106 ( .A(n2258), .Y(n4813) );
  BUFX2 U5107 ( .A(n2254), .Y(n4814) );
  BUFX2 U5108 ( .A(n2252), .Y(n4815) );
  BUFX2 U5109 ( .A(n2250), .Y(n4816) );
  BUFX2 U5110 ( .A(n2246), .Y(n4817) );
  BUFX2 U5111 ( .A(n2244), .Y(n4818) );
  BUFX2 U5112 ( .A(n2240), .Y(n4819) );
  BUFX2 U5113 ( .A(n11096), .Y(n4820) );
  BUFX2 U5114 ( .A(n11100), .Y(n4821) );
  BUFX2 U5115 ( .A(n11109), .Y(n4822) );
  BUFX2 U5116 ( .A(n11116), .Y(n4823) );
  BUFX2 U5117 ( .A(n11136), .Y(n4824) );
  BUFX2 U5118 ( .A(n11140), .Y(n4825) );
  BUFX2 U5119 ( .A(n11143), .Y(n4826) );
  BUFX2 U5120 ( .A(n11147), .Y(n4827) );
  BUFX2 U5121 ( .A(n11153), .Y(n4828) );
  BUFX2 U5122 ( .A(n11160), .Y(n4829) );
  BUFX2 U5123 ( .A(n11467), .Y(n4830) );
  BUFX2 U5124 ( .A(n11470), .Y(n4831) );
  BUFX2 U5125 ( .A(n11473), .Y(n4832) );
  BUFX2 U5126 ( .A(n11477), .Y(n4833) );
  BUFX2 U5127 ( .A(n11486), .Y(n4834) );
  BUFX2 U5128 ( .A(n11493), .Y(n4835) );
  BUFX2 U5129 ( .A(n11513), .Y(n4836) );
  BUFX2 U5130 ( .A(n11517), .Y(n4837) );
  BUFX2 U5131 ( .A(n11525), .Y(n4838) );
  BUFX2 U5132 ( .A(n11530), .Y(n4839) );
  BUFX2 U5133 ( .A(n11537), .Y(n4840) );
  BUFX2 U5134 ( .A(n11566), .Y(n4841) );
  BUFX2 U5135 ( .A(n11575), .Y(n4842) );
  BUFX2 U5136 ( .A(n11579), .Y(n4843) );
  BUFX2 U5137 ( .A(n11585), .Y(n4844) );
  BUFX2 U5138 ( .A(n11588), .Y(n4845) );
  BUFX2 U5139 ( .A(n11591), .Y(n4846) );
  BUFX2 U5140 ( .A(n11595), .Y(n4847) );
  BUFX2 U5141 ( .A(n11636), .Y(n4848) );
  BUFX2 U5142 ( .A(n11642), .Y(n4849) );
  BUFX2 U5143 ( .A(n11646), .Y(n4850) );
  BUFX2 U5144 ( .A(n11655), .Y(n4851) );
  BUFX2 U5145 ( .A(n11662), .Y(n4852) );
  BUFX2 U5146 ( .A(n11682), .Y(n4853) );
  BUFX2 U5147 ( .A(n11686), .Y(n4854) );
  BUFX2 U5148 ( .A(n11689), .Y(n4855) );
  BUFX2 U5149 ( .A(n11693), .Y(n4856) );
  BUFX2 U5150 ( .A(n11699), .Y(n4857) );
  BUFX2 U5151 ( .A(n11706), .Y(n4858) );
  BUFX2 U5152 ( .A(n11725), .Y(n4859) );
  BUFX2 U5153 ( .A(n11728), .Y(n4860) );
  BUFX2 U5154 ( .A(n11731), .Y(n4861) );
  BUFX2 U5155 ( .A(n11735), .Y(n4862) );
  BUFX2 U5156 ( .A(n11744), .Y(n4863) );
  BUFX2 U5157 ( .A(n11751), .Y(n4864) );
  BUFX2 U5158 ( .A(n11771), .Y(n4865) );
  BUFX2 U5159 ( .A(n11775), .Y(n4866) );
  BUFX2 U5160 ( .A(n11783), .Y(n4867) );
  BUFX2 U5161 ( .A(n11788), .Y(n4868) );
  BUFX2 U5162 ( .A(n11795), .Y(n4869) );
  BUFX2 U5163 ( .A(n11820), .Y(n4870) );
  BUFX2 U5164 ( .A(n11824), .Y(n4871) );
  BUFX2 U5165 ( .A(n11833), .Y(n4872) );
  BUFX2 U5166 ( .A(n11840), .Y(n4873) );
  BUFX2 U5167 ( .A(n11860), .Y(n4874) );
  BUFX2 U5168 ( .A(n11864), .Y(n4875) );
  BUFX2 U5169 ( .A(n11867), .Y(n4876) );
  BUFX2 U5170 ( .A(n11871), .Y(n4877) );
  BUFX2 U5171 ( .A(n11877), .Y(n4878) );
  BUFX2 U5172 ( .A(n11884), .Y(n4879) );
  BUFX2 U5173 ( .A(n11922), .Y(n4880) );
  BUFX2 U5174 ( .A(n11928), .Y(n4881) );
  BUFX2 U5175 ( .A(n11932), .Y(n4882) );
  BUFX2 U5176 ( .A(n11941), .Y(n4883) );
  BUFX2 U5177 ( .A(n11948), .Y(n4884) );
  BUFX2 U5178 ( .A(n11968), .Y(n4885) );
  BUFX2 U5179 ( .A(n11972), .Y(n4886) );
  BUFX2 U5180 ( .A(n11975), .Y(n4887) );
  BUFX2 U5181 ( .A(n11979), .Y(n4888) );
  BUFX2 U5182 ( .A(n11985), .Y(n4889) );
  BUFX2 U5183 ( .A(n11992), .Y(n4890) );
  BUFX2 U5184 ( .A(n12011), .Y(n4891) );
  BUFX2 U5185 ( .A(n12017), .Y(n4892) );
  BUFX2 U5186 ( .A(n12021), .Y(n4893) );
  BUFX2 U5187 ( .A(n12030), .Y(n4894) );
  BUFX2 U5188 ( .A(n12037), .Y(n4895) );
  BUFX2 U5189 ( .A(n12057), .Y(n4896) );
  BUFX2 U5190 ( .A(n12061), .Y(n4897) );
  BUFX2 U5191 ( .A(n12064), .Y(n4898) );
  BUFX2 U5192 ( .A(n12068), .Y(n4899) );
  BUFX2 U5193 ( .A(n12074), .Y(n4900) );
  BUFX2 U5194 ( .A(n12081), .Y(n4901) );
  BUFX2 U5195 ( .A(n12106), .Y(n4902) );
  BUFX2 U5196 ( .A(n12110), .Y(n4903) );
  BUFX2 U5197 ( .A(n12119), .Y(n4904) );
  BUFX2 U5198 ( .A(n12126), .Y(n4905) );
  BUFX2 U5199 ( .A(n12146), .Y(n4906) );
  BUFX2 U5200 ( .A(n12150), .Y(n4907) );
  BUFX2 U5201 ( .A(n12153), .Y(n4908) );
  BUFX2 U5202 ( .A(n12157), .Y(n4909) );
  BUFX2 U5203 ( .A(n12163), .Y(n4910) );
  BUFX2 U5204 ( .A(n12170), .Y(n4911) );
  BUFX2 U5205 ( .A(n12199), .Y(n4912) );
  BUFX2 U5206 ( .A(n12208), .Y(n4913) );
  BUFX2 U5207 ( .A(n12212), .Y(n4914) );
  BUFX2 U5208 ( .A(n12218), .Y(n4915) );
  BUFX2 U5209 ( .A(n12221), .Y(n4916) );
  BUFX2 U5210 ( .A(n12224), .Y(n4917) );
  BUFX2 U5211 ( .A(n12228), .Y(n4918) );
  BUFX2 U5212 ( .A(\Decision_AXILiteS_s_axi_U/n331 ), .Y(n4919) );
  BUFX2 U5213 ( .A(\Decision_AXILiteS_s_axi_U/n337 ), .Y(n4920) );
  BUFX2 U5214 ( .A(\Decision_AXILiteS_s_axi_U/n603 ), .Y(n4921) );
  BUFX2 U5215 ( .A(\Decision_AXILiteS_s_axi_U/n608 ), .Y(n4922) );
  BUFX2 U5216 ( .A(\Decision_AXILiteS_s_axi_U/n609 ), .Y(n4923) );
  BUFX2 U5217 ( .A(\Decision_AXILiteS_s_axi_U/n613 ), .Y(n4924) );
  BUFX2 U5218 ( .A(\Decision_AXILiteS_s_axi_U/n619 ), .Y(n4925) );
  BUFX2 U5219 ( .A(\Decision_AXILiteS_s_axi_U/n624 ), .Y(n4926) );
  AND2X1 U5220 ( .A(n5208), .B(n10514), .Y(n11169) );
  INVX1 U5221 ( .A(n11169), .Y(n4927) );
  AND2X1 U5222 ( .A(n5209), .B(n9740), .Y(n11546) );
  INVX1 U5223 ( .A(n11546), .Y(n4928) );
  AND2X1 U5224 ( .A(n9488), .B(n5942), .Y(n11626) );
  INVX1 U5225 ( .A(n11626), .Y(n4929) );
  AND2X1 U5226 ( .A(n5210), .B(n9622), .Y(n11715) );
  INVX1 U5227 ( .A(n11715), .Y(n4930) );
  AND2X1 U5228 ( .A(n5211), .B(n9322), .Y(n11804) );
  INVX1 U5229 ( .A(n11804), .Y(n4931) );
  AND2X1 U5230 ( .A(n5212), .B(n10430), .Y(n11893) );
  INVX1 U5231 ( .A(n11893), .Y(n4932) );
  AND2X1 U5232 ( .A(n5213), .B(n9623), .Y(n12001) );
  INVX1 U5233 ( .A(n12001), .Y(n4933) );
  AND2X1 U5234 ( .A(n5214), .B(n9736), .Y(n12090) );
  INVX1 U5235 ( .A(n12090), .Y(n4934) );
  AND2X1 U5236 ( .A(n5215), .B(n9737), .Y(n12179) );
  INVX1 U5237 ( .A(n12179), .Y(n4935) );
  AND2X1 U5238 ( .A(n9525), .B(n5945), .Y(n12259) );
  INVX1 U5239 ( .A(n12259), .Y(n4936) );
  AND2X1 U5240 ( .A(n10275), .B(n10274), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n13 ) );
  INVX1 U5241 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n13 ), 
        .Y(n4937) );
  AND2X1 U5242 ( .A(\recentVBools_data_q1[0] ), .B(n10056), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n3 ) );
  INVX1 U5243 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n3 ), 
        .Y(n4938) );
  AND2X1 U5244 ( .A(data[15]), .B(n8409), .Y(\Decision_AXILiteS_s_axi_U/n342 )
         );
  INVX1 U5245 ( .A(\Decision_AXILiteS_s_axi_U/n342 ), .Y(n4939) );
  AND2X1 U5246 ( .A(data[14]), .B(n8409), .Y(\Decision_AXILiteS_s_axi_U/n344 )
         );
  INVX1 U5247 ( .A(\Decision_AXILiteS_s_axi_U/n344 ), .Y(n4940) );
  AND2X1 U5248 ( .A(data[13]), .B(n8409), .Y(\Decision_AXILiteS_s_axi_U/n345 )
         );
  INVX1 U5249 ( .A(\Decision_AXILiteS_s_axi_U/n345 ), .Y(n4941) );
  AND2X1 U5250 ( .A(data[12]), .B(n8409), .Y(\Decision_AXILiteS_s_axi_U/n346 )
         );
  INVX1 U5251 ( .A(\Decision_AXILiteS_s_axi_U/n346 ), .Y(n4942) );
  AND2X1 U5252 ( .A(data[11]), .B(n8409), .Y(\Decision_AXILiteS_s_axi_U/n347 )
         );
  INVX1 U5253 ( .A(\Decision_AXILiteS_s_axi_U/n347 ), .Y(n4943) );
  AND2X1 U5254 ( .A(data[10]), .B(n8409), .Y(\Decision_AXILiteS_s_axi_U/n348 )
         );
  INVX1 U5255 ( .A(\Decision_AXILiteS_s_axi_U/n348 ), .Y(n4944) );
  AND2X1 U5256 ( .A(data[9]), .B(n8409), .Y(\Decision_AXILiteS_s_axi_U/n349 )
         );
  INVX1 U5257 ( .A(\Decision_AXILiteS_s_axi_U/n349 ), .Y(n4945) );
  AND2X1 U5258 ( .A(data[8]), .B(n8409), .Y(\Decision_AXILiteS_s_axi_U/n350 )
         );
  INVX1 U5259 ( .A(\Decision_AXILiteS_s_axi_U/n350 ), .Y(n4946) );
  AND2X1 U5260 ( .A(v_length[30]), .B(n8410), .Y(
        \Decision_AXILiteS_s_axi_U/n376 ) );
  INVX1 U5261 ( .A(\Decision_AXILiteS_s_axi_U/n376 ), .Y(n4947) );
  AND2X1 U5262 ( .A(v_length[28]), .B(n8410), .Y(
        \Decision_AXILiteS_s_axi_U/n378 ) );
  INVX1 U5263 ( .A(\Decision_AXILiteS_s_axi_U/n378 ), .Y(n4948) );
  AND2X1 U5264 ( .A(v_length[27]), .B(n8410), .Y(
        \Decision_AXILiteS_s_axi_U/n379 ) );
  INVX1 U5265 ( .A(\Decision_AXILiteS_s_axi_U/n379 ), .Y(n4949) );
  AND2X1 U5266 ( .A(v_length[26]), .B(n8410), .Y(
        \Decision_AXILiteS_s_axi_U/n380 ) );
  INVX1 U5267 ( .A(\Decision_AXILiteS_s_axi_U/n380 ), .Y(n4950) );
  AND2X1 U5268 ( .A(v_length[25]), .B(n8410), .Y(
        \Decision_AXILiteS_s_axi_U/n381 ) );
  INVX1 U5269 ( .A(\Decision_AXILiteS_s_axi_U/n381 ), .Y(n4951) );
  AND2X1 U5270 ( .A(v_length[24]), .B(n8410), .Y(
        \Decision_AXILiteS_s_axi_U/n382 ) );
  INVX1 U5271 ( .A(\Decision_AXILiteS_s_axi_U/n382 ), .Y(n4952) );
  AND2X1 U5272 ( .A(v_length[23]), .B(n6949), .Y(
        \Decision_AXILiteS_s_axi_U/n387 ) );
  INVX1 U5273 ( .A(\Decision_AXILiteS_s_axi_U/n387 ), .Y(n4953) );
  AND2X1 U5274 ( .A(v_length[22]), .B(n6949), .Y(
        \Decision_AXILiteS_s_axi_U/n389 ) );
  INVX1 U5275 ( .A(\Decision_AXILiteS_s_axi_U/n389 ), .Y(n4954) );
  AND2X1 U5276 ( .A(v_length[21]), .B(n6949), .Y(
        \Decision_AXILiteS_s_axi_U/n390 ) );
  INVX1 U5277 ( .A(\Decision_AXILiteS_s_axi_U/n390 ), .Y(n4955) );
  AND2X1 U5278 ( .A(v_length[20]), .B(n6949), .Y(
        \Decision_AXILiteS_s_axi_U/n391 ) );
  INVX1 U5279 ( .A(\Decision_AXILiteS_s_axi_U/n391 ), .Y(n4956) );
  AND2X1 U5280 ( .A(v_length[19]), .B(n6949), .Y(
        \Decision_AXILiteS_s_axi_U/n392 ) );
  INVX1 U5281 ( .A(\Decision_AXILiteS_s_axi_U/n392 ), .Y(n4957) );
  AND2X1 U5282 ( .A(v_length[18]), .B(n6949), .Y(
        \Decision_AXILiteS_s_axi_U/n393 ) );
  INVX1 U5283 ( .A(\Decision_AXILiteS_s_axi_U/n393 ), .Y(n4958) );
  AND2X1 U5284 ( .A(v_length[17]), .B(n6949), .Y(
        \Decision_AXILiteS_s_axi_U/n394 ) );
  INVX1 U5285 ( .A(\Decision_AXILiteS_s_axi_U/n394 ), .Y(n4959) );
  AND2X1 U5286 ( .A(v_length[16]), .B(n6949), .Y(
        \Decision_AXILiteS_s_axi_U/n395 ) );
  INVX1 U5287 ( .A(\Decision_AXILiteS_s_axi_U/n395 ), .Y(n4960) );
  AND2X1 U5288 ( .A(v_length[15]), .B(n7102), .Y(
        \Decision_AXILiteS_s_axi_U/n399 ) );
  INVX1 U5289 ( .A(\Decision_AXILiteS_s_axi_U/n399 ), .Y(n4961) );
  AND2X1 U5290 ( .A(v_length[14]), .B(n7102), .Y(
        \Decision_AXILiteS_s_axi_U/n401 ) );
  INVX1 U5291 ( .A(\Decision_AXILiteS_s_axi_U/n401 ), .Y(n4962) );
  AND2X1 U5292 ( .A(v_length[13]), .B(n7102), .Y(
        \Decision_AXILiteS_s_axi_U/n402 ) );
  INVX1 U5293 ( .A(\Decision_AXILiteS_s_axi_U/n402 ), .Y(n4963) );
  AND2X1 U5294 ( .A(v_length[12]), .B(n7102), .Y(
        \Decision_AXILiteS_s_axi_U/n403 ) );
  INVX1 U5295 ( .A(\Decision_AXILiteS_s_axi_U/n403 ), .Y(n4964) );
  AND2X1 U5296 ( .A(v_length[11]), .B(n7102), .Y(
        \Decision_AXILiteS_s_axi_U/n404 ) );
  INVX1 U5297 ( .A(\Decision_AXILiteS_s_axi_U/n404 ), .Y(n4965) );
  AND2X1 U5298 ( .A(v_length[10]), .B(n7102), .Y(
        \Decision_AXILiteS_s_axi_U/n405 ) );
  INVX1 U5299 ( .A(\Decision_AXILiteS_s_axi_U/n405 ), .Y(n4966) );
  AND2X1 U5300 ( .A(v_length[9]), .B(n7102), .Y(
        \Decision_AXILiteS_s_axi_U/n406 ) );
  INVX1 U5301 ( .A(\Decision_AXILiteS_s_axi_U/n406 ), .Y(n4967) );
  AND2X1 U5302 ( .A(v_length[8]), .B(n7102), .Y(
        \Decision_AXILiteS_s_axi_U/n407 ) );
  INVX1 U5303 ( .A(\Decision_AXILiteS_s_axi_U/n407 ), .Y(n4968) );
  AND2X1 U5304 ( .A(a_length[23]), .B(n7103), .Y(
        \Decision_AXILiteS_s_axi_U/n431 ) );
  INVX1 U5305 ( .A(\Decision_AXILiteS_s_axi_U/n431 ), .Y(n4969) );
  AND2X1 U5306 ( .A(a_length[22]), .B(n7103), .Y(
        \Decision_AXILiteS_s_axi_U/n433 ) );
  INVX1 U5307 ( .A(\Decision_AXILiteS_s_axi_U/n433 ), .Y(n4970) );
  AND2X1 U5308 ( .A(a_length[21]), .B(n7103), .Y(
        \Decision_AXILiteS_s_axi_U/n434 ) );
  INVX1 U5309 ( .A(\Decision_AXILiteS_s_axi_U/n434 ), .Y(n4971) );
  AND2X1 U5310 ( .A(a_length[20]), .B(n7103), .Y(
        \Decision_AXILiteS_s_axi_U/n435 ) );
  INVX1 U5311 ( .A(\Decision_AXILiteS_s_axi_U/n435 ), .Y(n4972) );
  AND2X1 U5312 ( .A(a_length[19]), .B(n7103), .Y(
        \Decision_AXILiteS_s_axi_U/n436 ) );
  INVX1 U5313 ( .A(\Decision_AXILiteS_s_axi_U/n436 ), .Y(n4973) );
  AND2X1 U5314 ( .A(a_length[18]), .B(n7103), .Y(
        \Decision_AXILiteS_s_axi_U/n437 ) );
  INVX1 U5315 ( .A(\Decision_AXILiteS_s_axi_U/n437 ), .Y(n4974) );
  AND2X1 U5316 ( .A(a_length[17]), .B(n7103), .Y(
        \Decision_AXILiteS_s_axi_U/n438 ) );
  INVX1 U5317 ( .A(\Decision_AXILiteS_s_axi_U/n438 ), .Y(n4975) );
  AND2X1 U5318 ( .A(a_length[16]), .B(n7103), .Y(
        \Decision_AXILiteS_s_axi_U/n439 ) );
  INVX1 U5319 ( .A(\Decision_AXILiteS_s_axi_U/n439 ), .Y(n4976) );
  AND2X1 U5320 ( .A(a_length[15]), .B(n6950), .Y(
        \Decision_AXILiteS_s_axi_U/n441 ) );
  INVX1 U5321 ( .A(\Decision_AXILiteS_s_axi_U/n441 ), .Y(n4977) );
  AND2X1 U5322 ( .A(a_length[14]), .B(n6950), .Y(
        \Decision_AXILiteS_s_axi_U/n443 ) );
  INVX1 U5323 ( .A(\Decision_AXILiteS_s_axi_U/n443 ), .Y(n4978) );
  AND2X1 U5324 ( .A(a_length[13]), .B(n6950), .Y(
        \Decision_AXILiteS_s_axi_U/n444 ) );
  INVX1 U5325 ( .A(\Decision_AXILiteS_s_axi_U/n444 ), .Y(n4979) );
  AND2X1 U5326 ( .A(a_length[12]), .B(n6950), .Y(
        \Decision_AXILiteS_s_axi_U/n445 ) );
  INVX1 U5327 ( .A(\Decision_AXILiteS_s_axi_U/n445 ), .Y(n4980) );
  AND2X1 U5328 ( .A(a_length[11]), .B(n6950), .Y(
        \Decision_AXILiteS_s_axi_U/n446 ) );
  INVX1 U5329 ( .A(\Decision_AXILiteS_s_axi_U/n446 ), .Y(n4981) );
  AND2X1 U5330 ( .A(a_length[10]), .B(n6950), .Y(
        \Decision_AXILiteS_s_axi_U/n447 ) );
  INVX1 U5331 ( .A(\Decision_AXILiteS_s_axi_U/n447 ), .Y(n4982) );
  AND2X1 U5332 ( .A(a_length[9]), .B(n6950), .Y(
        \Decision_AXILiteS_s_axi_U/n448 ) );
  INVX1 U5333 ( .A(\Decision_AXILiteS_s_axi_U/n448 ), .Y(n4983) );
  AND2X1 U5334 ( .A(a_length[8]), .B(n6950), .Y(
        \Decision_AXILiteS_s_axi_U/n449 ) );
  INVX1 U5335 ( .A(\Decision_AXILiteS_s_axi_U/n449 ), .Y(n4984) );
  AND2X1 U5336 ( .A(\Decision_AXILiteS_s_axi_U/n356 ), .B(
        \Decision_AXILiteS_s_axi_U/n473 ), .Y(\Decision_AXILiteS_s_axi_U/n472 ) );
  INVX1 U5337 ( .A(\Decision_AXILiteS_s_axi_U/n472 ), .Y(n4985) );
  AND2X1 U5338 ( .A(\Decision_AXILiteS_s_axi_U/n358 ), .B(
        \Decision_AXILiteS_s_axi_U/n473 ), .Y(\Decision_AXILiteS_s_axi_U/n474 ) );
  INVX1 U5339 ( .A(\Decision_AXILiteS_s_axi_U/n474 ), .Y(n4986) );
  AND2X1 U5340 ( .A(\Decision_AXILiteS_s_axi_U/n360 ), .B(
        \Decision_AXILiteS_s_axi_U/n473 ), .Y(\Decision_AXILiteS_s_axi_U/n475 ) );
  INVX1 U5341 ( .A(\Decision_AXILiteS_s_axi_U/n475 ), .Y(n4987) );
  AND2X1 U5342 ( .A(\Decision_AXILiteS_s_axi_U/n362 ), .B(
        \Decision_AXILiteS_s_axi_U/n473 ), .Y(\Decision_AXILiteS_s_axi_U/n476 ) );
  INVX1 U5343 ( .A(\Decision_AXILiteS_s_axi_U/n476 ), .Y(n4988) );
  AND2X1 U5344 ( .A(\Decision_AXILiteS_s_axi_U/n364 ), .B(
        \Decision_AXILiteS_s_axi_U/n473 ), .Y(\Decision_AXILiteS_s_axi_U/n477 ) );
  INVX1 U5345 ( .A(\Decision_AXILiteS_s_axi_U/n477 ), .Y(n4989) );
  AND2X1 U5346 ( .A(\Decision_AXILiteS_s_axi_U/n366 ), .B(
        \Decision_AXILiteS_s_axi_U/n473 ), .Y(\Decision_AXILiteS_s_axi_U/n478 ) );
  INVX1 U5347 ( .A(\Decision_AXILiteS_s_axi_U/n478 ), .Y(n4990) );
  AND2X1 U5348 ( .A(\Decision_AXILiteS_s_axi_U/n368 ), .B(
        \Decision_AXILiteS_s_axi_U/n473 ), .Y(\Decision_AXILiteS_s_axi_U/n479 ) );
  INVX1 U5349 ( .A(\Decision_AXILiteS_s_axi_U/n479 ), .Y(n4991) );
  AND2X1 U5350 ( .A(\Decision_AXILiteS_s_axi_U/n564 ), .B(
        \Decision_AXILiteS_s_axi_U/n473 ), .Y(\Decision_AXILiteS_s_axi_U/n480 ) );
  INVX1 U5351 ( .A(\Decision_AXILiteS_s_axi_U/n480 ), .Y(n4992) );
  AND2X1 U5352 ( .A(vthresh[23]), .B(n7268), .Y(
        \Decision_AXILiteS_s_axi_U/n494 ) );
  INVX1 U5353 ( .A(\Decision_AXILiteS_s_axi_U/n494 ), .Y(n4993) );
  AND2X1 U5354 ( .A(vthresh[22]), .B(n7268), .Y(
        \Decision_AXILiteS_s_axi_U/n496 ) );
  INVX1 U5355 ( .A(\Decision_AXILiteS_s_axi_U/n496 ), .Y(n4994) );
  AND2X1 U5356 ( .A(vthresh[21]), .B(n7268), .Y(
        \Decision_AXILiteS_s_axi_U/n497 ) );
  INVX1 U5357 ( .A(\Decision_AXILiteS_s_axi_U/n497 ), .Y(n4995) );
  AND2X1 U5358 ( .A(vthresh[20]), .B(n7268), .Y(
        \Decision_AXILiteS_s_axi_U/n498 ) );
  INVX1 U5359 ( .A(\Decision_AXILiteS_s_axi_U/n498 ), .Y(n4996) );
  AND2X1 U5360 ( .A(vthresh[19]), .B(n7268), .Y(
        \Decision_AXILiteS_s_axi_U/n499 ) );
  INVX1 U5361 ( .A(\Decision_AXILiteS_s_axi_U/n499 ), .Y(n4997) );
  AND2X1 U5362 ( .A(vthresh[18]), .B(n7268), .Y(
        \Decision_AXILiteS_s_axi_U/n500 ) );
  INVX1 U5363 ( .A(\Decision_AXILiteS_s_axi_U/n500 ), .Y(n4998) );
  AND2X1 U5364 ( .A(vthresh[17]), .B(n7268), .Y(
        \Decision_AXILiteS_s_axi_U/n501 ) );
  INVX1 U5365 ( .A(\Decision_AXILiteS_s_axi_U/n501 ), .Y(n4999) );
  AND2X1 U5366 ( .A(vthresh[16]), .B(n7268), .Y(
        \Decision_AXILiteS_s_axi_U/n502 ) );
  INVX1 U5367 ( .A(\Decision_AXILiteS_s_axi_U/n502 ), .Y(n5000) );
  AND2X1 U5368 ( .A(vthresh[15]), .B(n7445), .Y(
        \Decision_AXILiteS_s_axi_U/n504 ) );
  INVX1 U5369 ( .A(\Decision_AXILiteS_s_axi_U/n504 ), .Y(n5001) );
  AND2X1 U5370 ( .A(vthresh[14]), .B(n7445), .Y(
        \Decision_AXILiteS_s_axi_U/n506 ) );
  INVX1 U5371 ( .A(\Decision_AXILiteS_s_axi_U/n506 ), .Y(n5002) );
  AND2X1 U5372 ( .A(vthresh[13]), .B(n7445), .Y(
        \Decision_AXILiteS_s_axi_U/n507 ) );
  INVX1 U5373 ( .A(\Decision_AXILiteS_s_axi_U/n507 ), .Y(n5003) );
  AND2X1 U5374 ( .A(vthresh[12]), .B(n7445), .Y(
        \Decision_AXILiteS_s_axi_U/n508 ) );
  INVX1 U5375 ( .A(\Decision_AXILiteS_s_axi_U/n508 ), .Y(n5004) );
  AND2X1 U5376 ( .A(vthresh[11]), .B(n7445), .Y(
        \Decision_AXILiteS_s_axi_U/n509 ) );
  INVX1 U5377 ( .A(\Decision_AXILiteS_s_axi_U/n509 ), .Y(n5005) );
  AND2X1 U5378 ( .A(vthresh[10]), .B(n7445), .Y(
        \Decision_AXILiteS_s_axi_U/n510 ) );
  INVX1 U5379 ( .A(\Decision_AXILiteS_s_axi_U/n510 ), .Y(n5006) );
  AND2X1 U5380 ( .A(vthresh[9]), .B(n7445), .Y(
        \Decision_AXILiteS_s_axi_U/n511 ) );
  INVX1 U5381 ( .A(\Decision_AXILiteS_s_axi_U/n511 ), .Y(n5007) );
  AND2X1 U5382 ( .A(vthresh[8]), .B(n7445), .Y(
        \Decision_AXILiteS_s_axi_U/n512 ) );
  INVX1 U5383 ( .A(\Decision_AXILiteS_s_axi_U/n512 ), .Y(n5008) );
  AND2X1 U5384 ( .A(athresh[31]), .B(n7651), .Y(
        \Decision_AXILiteS_s_axi_U/n524 ) );
  INVX1 U5385 ( .A(\Decision_AXILiteS_s_axi_U/n524 ), .Y(n5009) );
  AND2X1 U5386 ( .A(athresh[30]), .B(n7651), .Y(
        \Decision_AXILiteS_s_axi_U/n526 ) );
  INVX1 U5387 ( .A(\Decision_AXILiteS_s_axi_U/n526 ), .Y(n5010) );
  AND2X1 U5388 ( .A(athresh[29]), .B(n7651), .Y(
        \Decision_AXILiteS_s_axi_U/n527 ) );
  INVX1 U5389 ( .A(\Decision_AXILiteS_s_axi_U/n527 ), .Y(n5011) );
  AND2X1 U5390 ( .A(athresh[28]), .B(n7651), .Y(
        \Decision_AXILiteS_s_axi_U/n528 ) );
  INVX1 U5391 ( .A(\Decision_AXILiteS_s_axi_U/n528 ), .Y(n5012) );
  AND2X1 U5392 ( .A(athresh[27]), .B(n7651), .Y(
        \Decision_AXILiteS_s_axi_U/n529 ) );
  INVX1 U5393 ( .A(\Decision_AXILiteS_s_axi_U/n529 ), .Y(n5013) );
  AND2X1 U5394 ( .A(athresh[26]), .B(n7651), .Y(
        \Decision_AXILiteS_s_axi_U/n530 ) );
  INVX1 U5395 ( .A(\Decision_AXILiteS_s_axi_U/n530 ), .Y(n5014) );
  AND2X1 U5396 ( .A(athresh[25]), .B(n7651), .Y(
        \Decision_AXILiteS_s_axi_U/n531 ) );
  INVX1 U5397 ( .A(\Decision_AXILiteS_s_axi_U/n531 ), .Y(n5015) );
  AND2X1 U5398 ( .A(athresh[24]), .B(n7651), .Y(
        \Decision_AXILiteS_s_axi_U/n532 ) );
  INVX1 U5399 ( .A(\Decision_AXILiteS_s_axi_U/n532 ), .Y(n5016) );
  AND2X1 U5400 ( .A(athresh[23]), .B(n7446), .Y(
        \Decision_AXILiteS_s_axi_U/n536 ) );
  INVX1 U5401 ( .A(\Decision_AXILiteS_s_axi_U/n536 ), .Y(n5017) );
  AND2X1 U5402 ( .A(athresh[22]), .B(n7446), .Y(
        \Decision_AXILiteS_s_axi_U/n538 ) );
  INVX1 U5403 ( .A(\Decision_AXILiteS_s_axi_U/n538 ), .Y(n5018) );
  AND2X1 U5404 ( .A(athresh[21]), .B(n7446), .Y(
        \Decision_AXILiteS_s_axi_U/n539 ) );
  INVX1 U5405 ( .A(\Decision_AXILiteS_s_axi_U/n539 ), .Y(n5019) );
  AND2X1 U5406 ( .A(athresh[20]), .B(n7446), .Y(
        \Decision_AXILiteS_s_axi_U/n540 ) );
  INVX1 U5407 ( .A(\Decision_AXILiteS_s_axi_U/n540 ), .Y(n5020) );
  AND2X1 U5408 ( .A(athresh[19]), .B(n7446), .Y(
        \Decision_AXILiteS_s_axi_U/n541 ) );
  INVX1 U5409 ( .A(\Decision_AXILiteS_s_axi_U/n541 ), .Y(n5021) );
  AND2X1 U5410 ( .A(athresh[18]), .B(n7446), .Y(
        \Decision_AXILiteS_s_axi_U/n542 ) );
  INVX1 U5411 ( .A(\Decision_AXILiteS_s_axi_U/n542 ), .Y(n5022) );
  AND2X1 U5412 ( .A(athresh[17]), .B(n7446), .Y(
        \Decision_AXILiteS_s_axi_U/n543 ) );
  INVX1 U5413 ( .A(\Decision_AXILiteS_s_axi_U/n543 ), .Y(n5023) );
  AND2X1 U5414 ( .A(athresh[16]), .B(n7446), .Y(
        \Decision_AXILiteS_s_axi_U/n544 ) );
  INVX1 U5415 ( .A(\Decision_AXILiteS_s_axi_U/n544 ), .Y(n5024) );
  AND2X1 U5416 ( .A(athresh[15]), .B(n7269), .Y(
        \Decision_AXILiteS_s_axi_U/n546 ) );
  INVX1 U5417 ( .A(\Decision_AXILiteS_s_axi_U/n546 ), .Y(n5025) );
  AND2X1 U5418 ( .A(athresh[14]), .B(n7269), .Y(
        \Decision_AXILiteS_s_axi_U/n548 ) );
  INVX1 U5419 ( .A(\Decision_AXILiteS_s_axi_U/n548 ), .Y(n5026) );
  AND2X1 U5420 ( .A(athresh[13]), .B(n7269), .Y(
        \Decision_AXILiteS_s_axi_U/n549 ) );
  INVX1 U5421 ( .A(\Decision_AXILiteS_s_axi_U/n549 ), .Y(n5027) );
  AND2X1 U5422 ( .A(athresh[12]), .B(n7269), .Y(
        \Decision_AXILiteS_s_axi_U/n550 ) );
  INVX1 U5423 ( .A(\Decision_AXILiteS_s_axi_U/n550 ), .Y(n5028) );
  AND2X1 U5424 ( .A(athresh[11]), .B(n7269), .Y(
        \Decision_AXILiteS_s_axi_U/n551 ) );
  INVX1 U5425 ( .A(\Decision_AXILiteS_s_axi_U/n551 ), .Y(n5029) );
  AND2X1 U5426 ( .A(athresh[10]), .B(n7269), .Y(
        \Decision_AXILiteS_s_axi_U/n552 ) );
  INVX1 U5427 ( .A(\Decision_AXILiteS_s_axi_U/n552 ), .Y(n5030) );
  AND2X1 U5428 ( .A(athresh[9]), .B(n7269), .Y(
        \Decision_AXILiteS_s_axi_U/n553 ) );
  INVX1 U5429 ( .A(\Decision_AXILiteS_s_axi_U/n553 ), .Y(n5031) );
  AND2X1 U5430 ( .A(athresh[8]), .B(n7269), .Y(
        \Decision_AXILiteS_s_axi_U/n554 ) );
  INVX1 U5431 ( .A(\Decision_AXILiteS_s_axi_U/n554 ), .Y(n5032) );
  AND2X1 U5432 ( .A(n5948), .B(\Decision_AXILiteS_s_axi_U/n579 ), .Y(
        \Decision_AXILiteS_s_axi_U/n582 ) );
  INVX1 U5433 ( .A(\Decision_AXILiteS_s_axi_U/n582 ), .Y(n5033) );
  AND2X1 U5434 ( .A(n685), .B(\Decision_AXILiteS_s_axi_U/n579 ), .Y(
        \Decision_AXILiteS_s_axi_U/n590 ) );
  INVX1 U5435 ( .A(\Decision_AXILiteS_s_axi_U/n590 ), .Y(n5034) );
  AND2X1 U5436 ( .A(toReturn_1_fu_1395_p3_12), .B(
        \Decision_AXILiteS_s_axi_U/n579 ), .Y(\Decision_AXILiteS_s_axi_U/n594 ) );
  INVX1 U5437 ( .A(\Decision_AXILiteS_s_axi_U/n594 ), .Y(n5035) );
  AND2X1 U5438 ( .A(tmp_29_i1_fu_1065_p2[25]), .B(n8922), .Y(n3219) );
  INVX1 U5439 ( .A(n3219), .Y(n5036) );
  AND2X1 U5440 ( .A(tmp_29_i1_fu_1065_p2[26]), .B(n8922), .Y(n3218) );
  INVX1 U5441 ( .A(n3218), .Y(n5037) );
  AND2X1 U5442 ( .A(tmp_29_i1_fu_1065_p2[29]), .B(n8922), .Y(n3215) );
  INVX1 U5443 ( .A(n3215), .Y(n5038) );
  AND2X1 U5444 ( .A(tmp_29_i_fu_752_p2[25]), .B(n8920), .Y(n3167) );
  INVX1 U5445 ( .A(n3167), .Y(n5039) );
  AND2X1 U5446 ( .A(tmp_29_i_fu_752_p2[26]), .B(n8920), .Y(n3166) );
  INVX1 U5447 ( .A(n3166), .Y(n5040) );
  AND2X1 U5448 ( .A(tmp_29_i_fu_752_p2[29]), .B(n8920), .Y(n3163) );
  INVX1 U5449 ( .A(n3163), .Y(n5041) );
  AND2X1 U5450 ( .A(a_flip[3]), .B(n8952), .Y(n3145) );
  INVX1 U5451 ( .A(n3145), .Y(n5042) );
  AND2X1 U5452 ( .A(a_flip[4]), .B(n8951), .Y(n3144) );
  INVX1 U5453 ( .A(n3144), .Y(n5043) );
  AND2X1 U5454 ( .A(a_flip[6]), .B(n8951), .Y(n3140) );
  INVX1 U5455 ( .A(n3140), .Y(n5044) );
  AND2X1 U5456 ( .A(v_flip[2]), .B(n8952), .Y(n3134) );
  INVX1 U5457 ( .A(n3134), .Y(n5045) );
  AND2X1 U5458 ( .A(v_flip[3]), .B(n8952), .Y(n3133) );
  INVX1 U5459 ( .A(n3133), .Y(n5046) );
  AND2X1 U5460 ( .A(a_length[15]), .B(n8953), .Y(n3096) );
  INVX1 U5461 ( .A(n3096), .Y(n5047) );
  AND2X1 U5462 ( .A(a_length[16]), .B(n8953), .Y(n3094) );
  INVX1 U5463 ( .A(n3094), .Y(n5048) );
  AND2X1 U5464 ( .A(a_length[30]), .B(n8954), .Y(n3066) );
  INVX1 U5465 ( .A(n3066), .Y(n5049) );
  AND2X1 U5466 ( .A(a_length[31]), .B(n8954), .Y(n3064) );
  INVX1 U5467 ( .A(n3064), .Y(n5050) );
  AND2X1 U5468 ( .A(sum_reg_308[19]), .B(n8929), .Y(n2622) );
  INVX1 U5469 ( .A(n2622), .Y(n5051) );
  AND2X1 U5470 ( .A(sum_1_reg_376[19]), .B(n8930), .Y(n2484) );
  INVX1 U5471 ( .A(n2484), .Y(n5052) );
  AND2X1 U5472 ( .A(sum_1_reg_376[11]), .B(n8930), .Y(n2452) );
  INVX1 U5473 ( .A(n2452), .Y(n5053) );
  AND2X1 U5474 ( .A(recentdatapoints_head_i[6]), .B(n8977), .Y(n1977) );
  INVX1 U5475 ( .A(n1977), .Y(n5054) );
  AND2X1 U5476 ( .A(recentdatapoints_head_i[11]), .B(n8980), .Y(n1972) );
  INVX1 U5477 ( .A(n1972), .Y(n5055) );
  AND2X1 U5478 ( .A(recentdatapoints_head_i[18]), .B(n8979), .Y(n1965) );
  INVX1 U5479 ( .A(n1965), .Y(n5056) );
  AND2X1 U5480 ( .A(CircularBuffer_head_i_read_ass_reg_1624[0]), .B(n9011), 
        .Y(n1796) );
  INVX1 U5481 ( .A(n1796), .Y(n5057) );
  AND2X1 U5482 ( .A(n10024), .B(n8993), .Y(n1794) );
  INVX1 U5483 ( .A(n1794), .Y(n5058) );
  AND2X1 U5484 ( .A(CircularBuffer_head_i_read_ass_reg_1624[5]), .B(n9011), 
        .Y(n1790) );
  INVX1 U5485 ( .A(n1790), .Y(n5059) );
  AND2X1 U5486 ( .A(recentVBools_head_i[11]), .B(n9007), .Y(n1771) );
  INVX1 U5487 ( .A(n1771), .Y(n5060) );
  AND2X1 U5488 ( .A(CircularBuffer_head_i_read_ass_reg_1624[12]), .B(n9010), 
        .Y(n1769) );
  INVX1 U5489 ( .A(n1769), .Y(n5061) );
  AND2X1 U5490 ( .A(CircularBuffer_head_i_read_ass_reg_1624[27]), .B(n9008), 
        .Y(n1724) );
  INVX1 U5491 ( .A(n1724), .Y(n5062) );
  AND2X1 U5492 ( .A(recentVBools_head_i[27]), .B(n9008), .Y(n1723) );
  INVX1 U5493 ( .A(n1723), .Y(n5063) );
  AND2X1 U5494 ( .A(CircularBuffer_head_i_read_ass_reg_1624[28]), .B(n9008), 
        .Y(n1721) );
  INVX1 U5495 ( .A(n1721), .Y(n5064) );
  AND2X1 U5496 ( .A(\tmp_i3_reg_1674[0] ), .B(n9013), .Y(n1651) );
  INVX1 U5497 ( .A(n1651), .Y(n5065) );
  AND2X1 U5498 ( .A(n8991), .B(CircularBuffer_len_read_assign_1_fu_778_p3[1]), 
        .Y(n1644) );
  INVX1 U5499 ( .A(n1644), .Y(n5066) );
  AND2X1 U5500 ( .A(n8991), .B(CircularBuffer_len_read_assign_1_fu_778_p3[3]), 
        .Y(n1642) );
  INVX1 U5501 ( .A(n1642), .Y(n5067) );
  AND2X1 U5502 ( .A(n2784), .B(n8992), .Y(n1640) );
  INVX1 U5503 ( .A(n1640), .Y(n5068) );
  AND2X1 U5504 ( .A(n2776), .B(n8993), .Y(n1635) );
  INVX1 U5505 ( .A(n1635), .Y(n5069) );
  AND2X1 U5506 ( .A(n2754), .B(n8992), .Y(n1620) );
  INVX1 U5507 ( .A(n1620), .Y(n5070) );
  AND2X1 U5508 ( .A(n2752), .B(n8993), .Y(n1619) );
  INVX1 U5509 ( .A(n1619), .Y(n5071) );
  AND2X1 U5510 ( .A(n2750), .B(n8991), .Y(n1618) );
  INVX1 U5511 ( .A(n1618), .Y(n5072) );
  AND2X1 U5512 ( .A(n2746), .B(n8992), .Y(n1614) );
  INVX1 U5513 ( .A(n1614), .Y(n5073) );
  AND2X1 U5514 ( .A(n2738), .B(n8991), .Y(n1608) );
  INVX1 U5515 ( .A(n1608), .Y(n5074) );
  AND2X1 U5516 ( .A(n2736), .B(n8992), .Y(n1606) );
  INVX1 U5517 ( .A(n1606), .Y(n5075) );
  AND2X1 U5518 ( .A(CircularBuffer_len_write_assig_fu_817_p2[6]), .B(n8894), 
        .Y(n1594) );
  INVX1 U5519 ( .A(n1594), .Y(n5076) );
  AND2X1 U5520 ( .A(CircularBuffer_len_write_assig_fu_817_p2[12]), .B(n8894), 
        .Y(n1585) );
  INVX1 U5521 ( .A(n1585), .Y(n5077) );
  AND2X1 U5522 ( .A(CircularBuffer_len_write_assig_fu_817_p2[13]), .B(n8894), 
        .Y(n1583) );
  INVX1 U5523 ( .A(n1583), .Y(n5078) );
  AND2X1 U5524 ( .A(CircularBuffer_len_write_assig_fu_817_p2[16]), .B(n8894), 
        .Y(n1579) );
  INVX1 U5525 ( .A(n1579), .Y(n5079) );
  AND2X1 U5526 ( .A(CircularBuffer_len_write_assig_fu_817_p2[17]), .B(n8894), 
        .Y(n1578) );
  INVX1 U5527 ( .A(n1578), .Y(n5080) );
  AND2X1 U5528 ( .A(CircularBuffer_len_write_assig_fu_817_p2[18]), .B(n1646), 
        .Y(n1577) );
  INVX1 U5529 ( .A(n1577), .Y(n5081) );
  AND2X1 U5530 ( .A(CircularBuffer_len_write_assig_fu_817_p2[19]), .B(n8894), 
        .Y(n1575) );
  INVX1 U5531 ( .A(n1575), .Y(n5082) );
  AND2X1 U5532 ( .A(CircularBuffer_len_write_assig_fu_817_p2[20]), .B(n8894), 
        .Y(n1573) );
  INVX1 U5533 ( .A(n1573), .Y(n5083) );
  AND2X1 U5534 ( .A(CircularBuffer_len_write_assig_fu_817_p2[21]), .B(n1646), 
        .Y(n1572) );
  INVX1 U5535 ( .A(n1572), .Y(n5084) );
  AND2X1 U5536 ( .A(CircularBuffer_len_write_assig_fu_817_p2[22]), .B(n8894), 
        .Y(n1570) );
  INVX1 U5537 ( .A(n1570), .Y(n5085) );
  AND2X1 U5538 ( .A(CircularBuffer_len_write_assig_fu_817_p2[24]), .B(n8894), 
        .Y(n1567) );
  INVX1 U5539 ( .A(n1567), .Y(n5086) );
  AND2X1 U5540 ( .A(CircularBuffer_len_write_assig_fu_817_p2[25]), .B(n8894), 
        .Y(n1566) );
  INVX1 U5541 ( .A(n1566), .Y(n5087) );
  AND2X1 U5542 ( .A(CircularBuffer_len_write_assig_fu_817_p2[26]), .B(n8894), 
        .Y(n1564) );
  INVX1 U5543 ( .A(n1564), .Y(n5088) );
  AND2X1 U5544 ( .A(CircularBuffer_len_write_assig_fu_817_p2[27]), .B(n8894), 
        .Y(n1562) );
  INVX1 U5545 ( .A(n1562), .Y(n5089) );
  AND2X1 U5546 ( .A(CircularBuffer_len_write_assig_fu_817_p2[28]), .B(n1646), 
        .Y(n1561) );
  INVX1 U5547 ( .A(n1561), .Y(n5090) );
  AND2X1 U5548 ( .A(CircularBuffer_len_write_assig_fu_817_p2[29]), .B(n8894), 
        .Y(n1560) );
  INVX1 U5549 ( .A(n1560), .Y(n5091) );
  AND2X1 U5550 ( .A(CircularBuffer_len_write_assig_fu_817_p2[31]), .B(n1646), 
        .Y(n1556) );
  INVX1 U5551 ( .A(n1556), .Y(n5092) );
  AND2X1 U5552 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[30]), .B(n9034), 
        .Y(n1400) );
  INVX1 U5553 ( .A(n1400), .Y(n5093) );
  AND2X1 U5554 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[29]), .B(n9034), 
        .Y(n1398) );
  INVX1 U5555 ( .A(n1398), .Y(n5094) );
  AND2X1 U5556 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[27]), .B(n9032), 
        .Y(n1394) );
  INVX1 U5557 ( .A(n1394), .Y(n5095) );
  AND2X1 U5558 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[22]), .B(n9032), 
        .Y(n1384) );
  INVX1 U5559 ( .A(n1384), .Y(n5096) );
  AND2X1 U5560 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[21]), .B(n9032), 
        .Y(n1382) );
  INVX1 U5561 ( .A(n1382), .Y(n5097) );
  AND2X1 U5562 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[19]), .B(n9032), 
        .Y(n1378) );
  INVX1 U5563 ( .A(n1378), .Y(n5098) );
  AND2X1 U5564 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[17]), .B(n9033), 
        .Y(n1374) );
  INVX1 U5565 ( .A(n1374), .Y(n5099) );
  AND2X1 U5566 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[16]), .B(n9033), 
        .Y(n1372) );
  INVX1 U5567 ( .A(n1372), .Y(n5100) );
  AND2X1 U5568 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[15]), .B(n9033), 
        .Y(n1370) );
  INVX1 U5569 ( .A(n1370), .Y(n5101) );
  AND2X1 U5570 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[14]), .B(n9034), 
        .Y(n1368) );
  INVX1 U5571 ( .A(n1368), .Y(n5102) );
  AND2X1 U5572 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[13]), .B(n9034), 
        .Y(n1366) );
  INVX1 U5573 ( .A(n1366), .Y(n5103) );
  AND2X1 U5574 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[10]), .B(n9035), 
        .Y(n1360) );
  INVX1 U5575 ( .A(n1360), .Y(n5104) );
  AND2X1 U5576 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[9]), .B(n9035), 
        .Y(n1358) );
  INVX1 U5577 ( .A(n1358), .Y(n5105) );
  AND2X1 U5578 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[5]), .B(n9036), 
        .Y(n1350) );
  INVX1 U5579 ( .A(n1350), .Y(n5106) );
  AND2X1 U5580 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[5]), .B(n9037), 
        .Y(n1332) );
  INVX1 U5581 ( .A(n1332), .Y(n5107) );
  AND2X1 U5582 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[6]), .B(n9038), 
        .Y(n1330) );
  INVX1 U5583 ( .A(n1330), .Y(n5108) );
  AND2X1 U5584 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[9]), .B(n9039), 
        .Y(n1323) );
  INVX1 U5585 ( .A(n1323), .Y(n5109) );
  AND2X1 U5586 ( .A(tmp_5_fu_726_p2[18]), .B(n8994), .Y(n1136) );
  INVX1 U5587 ( .A(n1136), .Y(n5110) );
  AND2X1 U5588 ( .A(tmp_5_fu_726_p2[19]), .B(n8994), .Y(n1132) );
  INVX1 U5589 ( .A(n1132), .Y(n5111) );
  AND2X1 U5590 ( .A(tmp_5_fu_726_p2[20]), .B(n8994), .Y(n1128) );
  INVX1 U5591 ( .A(n1128), .Y(n5112) );
  AND2X1 U5592 ( .A(tmp_4_fu_716_p2[5]), .B(n8995), .Y(n1062) );
  INVX1 U5593 ( .A(n1062), .Y(n5113) );
  AND2X1 U5594 ( .A(tmp_4_fu_716_p2[6]), .B(n8995), .Y(n1059) );
  INVX1 U5595 ( .A(n1059), .Y(n5114) );
  AND2X1 U5596 ( .A(tmp_4_fu_716_p2[7]), .B(n8995), .Y(n1056) );
  INVX1 U5597 ( .A(n1056), .Y(n5115) );
  AND2X1 U5598 ( .A(tmp_4_fu_716_p2[24]), .B(n8996), .Y(n999) );
  INVX1 U5599 ( .A(n999), .Y(n5116) );
  AND2X1 U5600 ( .A(tmp_4_fu_716_p2[25]), .B(n8996), .Y(n995) );
  INVX1 U5601 ( .A(n995), .Y(n5117) );
  AND2X1 U5602 ( .A(tmp_4_fu_716_p2[26]), .B(n8996), .Y(n992) );
  INVX1 U5603 ( .A(n992), .Y(n5118) );
  AND2X1 U5604 ( .A(n2291), .B(n9018), .Y(n964) );
  INVX1 U5605 ( .A(n964), .Y(n5119) );
  AND2X1 U5606 ( .A(n2289), .B(n9018), .Y(n963) );
  INVX1 U5607 ( .A(n963), .Y(n5120) );
  AND2X1 U5608 ( .A(n2277), .B(n9018), .Y(n954) );
  INVX1 U5609 ( .A(n954), .Y(n5121) );
  AND2X1 U5610 ( .A(n2275), .B(n9018), .Y(n953) );
  INVX1 U5611 ( .A(n953), .Y(n5122) );
  AND2X1 U5612 ( .A(n2269), .B(n9017), .Y(n948) );
  INVX1 U5613 ( .A(n948), .Y(n5123) );
  AND2X1 U5614 ( .A(n2267), .B(n9017), .Y(n947) );
  INVX1 U5615 ( .A(n947), .Y(n5124) );
  AND2X1 U5616 ( .A(n2265), .B(n9018), .Y(n946) );
  INVX1 U5617 ( .A(n946), .Y(n5125) );
  AND2X1 U5618 ( .A(n2263), .B(n9018), .Y(n945) );
  INVX1 U5619 ( .A(n945), .Y(n5126) );
  AND2X1 U5620 ( .A(n2261), .B(n9018), .Y(n944) );
  INVX1 U5621 ( .A(n944), .Y(n5127) );
  AND2X1 U5622 ( .A(n2259), .B(n9018), .Y(n943) );
  INVX1 U5623 ( .A(n943), .Y(n5128) );
  AND2X1 U5624 ( .A(n2253), .B(n9018), .Y(n938) );
  INVX1 U5625 ( .A(n938), .Y(n5129) );
  AND2X1 U5626 ( .A(n2251), .B(n9018), .Y(n936) );
  INVX1 U5627 ( .A(n936), .Y(n5130) );
  AND2X1 U5628 ( .A(n2249), .B(n9018), .Y(n934) );
  INVX1 U5629 ( .A(n934), .Y(n5131) );
  AND2X1 U5630 ( .A(n2245), .B(n9018), .Y(n932) );
  INVX1 U5631 ( .A(n932), .Y(n5132) );
  AND2X1 U5632 ( .A(n2243), .B(n9018), .Y(n930) );
  INVX1 U5633 ( .A(n930), .Y(n5133) );
  AND2X1 U5634 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[6]), .B(n8891), 
        .Y(n918) );
  INVX1 U5635 ( .A(n918), .Y(n5134) );
  AND2X1 U5636 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[12]), .B(n8891), .Y(n909) );
  INVX1 U5637 ( .A(n909), .Y(n5135) );
  AND2X1 U5638 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[13]), .B(n8891), .Y(n907) );
  INVX1 U5639 ( .A(n907), .Y(n5136) );
  AND2X1 U5640 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[16]), .B(n8891), .Y(n903) );
  INVX1 U5641 ( .A(n903), .Y(n5137) );
  AND2X1 U5642 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[17]), .B(n8891), .Y(n902) );
  INVX1 U5643 ( .A(n902), .Y(n5138) );
  AND2X1 U5644 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[18]), .B(n970), 
        .Y(n901) );
  INVX1 U5645 ( .A(n901), .Y(n5139) );
  AND2X1 U5646 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[19]), .B(n8891), .Y(n899) );
  INVX1 U5647 ( .A(n899), .Y(n5140) );
  AND2X1 U5648 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[20]), .B(n8891), .Y(n897) );
  INVX1 U5649 ( .A(n897), .Y(n5141) );
  AND2X1 U5650 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[21]), .B(n970), 
        .Y(n896) );
  INVX1 U5651 ( .A(n896), .Y(n5142) );
  AND2X1 U5652 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[22]), .B(n8891), .Y(n894) );
  INVX1 U5653 ( .A(n894), .Y(n5143) );
  AND2X1 U5654 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[24]), .B(n8891), .Y(n891) );
  INVX1 U5655 ( .A(n891), .Y(n5144) );
  AND2X1 U5656 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[25]), .B(n8891), .Y(n890) );
  INVX1 U5657 ( .A(n890), .Y(n5145) );
  AND2X1 U5658 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[26]), .B(n8891), .Y(n888) );
  INVX1 U5659 ( .A(n888), .Y(n5146) );
  AND2X1 U5660 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[27]), .B(n8891), .Y(n886) );
  INVX1 U5661 ( .A(n886), .Y(n5147) );
  AND2X1 U5662 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[28]), .B(n970), 
        .Y(n885) );
  INVX1 U5663 ( .A(n885), .Y(n5148) );
  AND2X1 U5664 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[29]), .B(n8891), .Y(n884) );
  INVX1 U5665 ( .A(n884), .Y(n5149) );
  AND2X1 U5666 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[31]), .B(n970), 
        .Y(n880) );
  INVX1 U5667 ( .A(n880), .Y(n5150) );
  AND2X1 U5668 ( .A(AbeatDelay[0]), .B(n8896), .Y(n793) );
  INVX1 U5669 ( .A(n793), .Y(n5151) );
  AND2X1 U5670 ( .A(AbeatDelay[4]), .B(n8896), .Y(n777) );
  INVX1 U5671 ( .A(n777), .Y(n5152) );
  AND2X1 U5672 ( .A(tmp_3_fu_706_p2[11]), .B(n8997), .Y(n757) );
  INVX1 U5673 ( .A(n757), .Y(n5153) );
  AND2X1 U5674 ( .A(tmp_3_fu_706_p2[12]), .B(n8997), .Y(n753) );
  INVX1 U5675 ( .A(n753), .Y(n5154) );
  AND2X1 U5676 ( .A(AbeatDelay[12]), .B(n10670), .Y(n751) );
  INVX1 U5677 ( .A(n751), .Y(n5155) );
  AND2X1 U5678 ( .A(tmp_3_fu_706_p2[13]), .B(n8997), .Y(n749) );
  INVX1 U5679 ( .A(n749), .Y(n5156) );
  AND2X1 U5680 ( .A(AstimDelay[6]), .B(n8896), .Y(n665) );
  INVX1 U5681 ( .A(n665), .Y(n5157) );
  AND2X1 U5682 ( .A(tmp_6_fu_497_p3[9]), .B(n8966), .Y(n657) );
  INVX1 U5683 ( .A(n657), .Y(n5158) );
  AND2X1 U5684 ( .A(tmp_6_fu_497_p3[10]), .B(n8966), .Y(n654) );
  INVX1 U5685 ( .A(n654), .Y(n5159) );
  AND2X1 U5686 ( .A(AstimDelay[23]), .B(n8896), .Y(n614) );
  INVX1 U5687 ( .A(n614), .Y(n5160) );
  AND2X1 U5688 ( .A(tmp_6_fu_497_p3[27]), .B(n8965), .Y(n603) );
  INVX1 U5689 ( .A(n603), .Y(n5161) );
  AND2X1 U5690 ( .A(tmp_6_fu_497_p3[28]), .B(n8965), .Y(n600) );
  INVX1 U5691 ( .A(n600), .Y(n5162) );
  AND2X1 U5692 ( .A(tmp_6_fu_497_p3[29]), .B(n8965), .Y(n597) );
  INVX1 U5693 ( .A(n597), .Y(n5163) );
  AND2X1 U5694 ( .A(tmp_6_fu_497_p3[30]), .B(n8965), .Y(n594) );
  INVX1 U5695 ( .A(n594), .Y(n5164) );
  AND2X1 U5696 ( .A(n10776), .B(n8965), .Y(n583) );
  INVX1 U5697 ( .A(n583), .Y(n5165) );
  AND2X1 U5698 ( .A(VstimDelay[9]), .B(n8896), .Y(n556) );
  INVX1 U5699 ( .A(n556), .Y(n5166) );
  AND2X1 U5700 ( .A(tmp_7_fu_511_p3[11]), .B(n8964), .Y(n551) );
  INVX1 U5701 ( .A(n551), .Y(n5167) );
  AND2X1 U5702 ( .A(tmp_7_fu_511_p3[12]), .B(n8964), .Y(n548) );
  INVX1 U5703 ( .A(n548), .Y(n5168) );
  AND2X1 U5704 ( .A(datapointA_1_fu_1017_p2[10]), .B(n439), .Y(n470) );
  INVX1 U5705 ( .A(n470), .Y(n5169) );
  AND2X1 U5706 ( .A(datapointA_1_fu_1017_p2[11]), .B(n439), .Y(n468) );
  INVX1 U5707 ( .A(n468), .Y(n5170) );
  AND2X1 U5708 ( .A(datapointA_1_fu_1017_p2[12]), .B(n439), .Y(n466) );
  INVX1 U5709 ( .A(n466), .Y(n5171) );
  AND2X1 U5710 ( .A(datapointA_1_fu_1017_p2[13]), .B(n439), .Y(n464) );
  INVX1 U5711 ( .A(n464), .Y(n5172) );
  AND2X1 U5712 ( .A(datapointA_1_fu_1017_p2[14]), .B(n439), .Y(n462) );
  INVX1 U5713 ( .A(n462), .Y(n5173) );
  AND2X1 U5714 ( .A(datapointA_1_fu_1017_p2[15]), .B(n439), .Y(n460) );
  INVX1 U5715 ( .A(n460), .Y(n5174) );
  AND2X1 U5716 ( .A(datapointA_1_fu_1017_p2[1]), .B(n439), .Y(n459) );
  INVX1 U5717 ( .A(n459), .Y(n5175) );
  AND2X1 U5718 ( .A(datapointA_1_fu_1017_p2[2]), .B(n439), .Y(n457) );
  INVX1 U5719 ( .A(n457), .Y(n5176) );
  AND2X1 U5720 ( .A(datapointA_1_fu_1017_p2[3]), .B(n439), .Y(n455) );
  INVX1 U5721 ( .A(n455), .Y(n5177) );
  AND2X1 U5722 ( .A(datapointA_1_fu_1017_p2[4]), .B(n439), .Y(n453) );
  INVX1 U5723 ( .A(n453), .Y(n5178) );
  AND2X1 U5724 ( .A(datapointA_1_fu_1017_p2[5]), .B(n439), .Y(n451) );
  INVX1 U5725 ( .A(n451), .Y(n5179) );
  AND2X1 U5726 ( .A(datapointA_1_fu_1017_p2[6]), .B(n439), .Y(n449) );
  INVX1 U5727 ( .A(n449), .Y(n5180) );
  AND2X1 U5728 ( .A(datapointA_1_fu_1017_p2[7]), .B(n439), .Y(n447) );
  INVX1 U5729 ( .A(n447), .Y(n5181) );
  AND2X1 U5730 ( .A(datapointA_1_fu_1017_p2[8]), .B(n439), .Y(n445) );
  INVX1 U5731 ( .A(n445), .Y(n5182) );
  AND2X1 U5732 ( .A(datapointA_1_fu_1017_p2[9]), .B(n439), .Y(n443) );
  INVX1 U5733 ( .A(n443), .Y(n5183) );
  AND2X1 U5734 ( .A(datapointV_1_fu_674_p2[10]), .B(n397), .Y(n428) );
  INVX1 U5735 ( .A(n428), .Y(n5184) );
  AND2X1 U5736 ( .A(datapointV_1_fu_674_p2[11]), .B(n397), .Y(n426) );
  INVX1 U5737 ( .A(n426), .Y(n5185) );
  AND2X1 U5738 ( .A(datapointV_1_fu_674_p2[12]), .B(n397), .Y(n424) );
  INVX1 U5739 ( .A(n424), .Y(n5186) );
  AND2X1 U5740 ( .A(datapointV_1_fu_674_p2[13]), .B(n397), .Y(n422) );
  INVX1 U5741 ( .A(n422), .Y(n5187) );
  AND2X1 U5742 ( .A(datapointV_1_fu_674_p2[14]), .B(n397), .Y(n420) );
  INVX1 U5743 ( .A(n420), .Y(n5188) );
  AND2X1 U5744 ( .A(datapointV_1_fu_674_p2[15]), .B(n397), .Y(n418) );
  INVX1 U5745 ( .A(n418), .Y(n5189) );
  AND2X1 U5746 ( .A(datapointV_1_fu_674_p2[1]), .B(n397), .Y(n417) );
  INVX1 U5747 ( .A(n417), .Y(n5190) );
  AND2X1 U5748 ( .A(datapointV_1_fu_674_p2[2]), .B(n397), .Y(n415) );
  INVX1 U5749 ( .A(n415), .Y(n5191) );
  AND2X1 U5750 ( .A(datapointV_1_fu_674_p2[3]), .B(n397), .Y(n413) );
  INVX1 U5751 ( .A(n413), .Y(n5192) );
  AND2X1 U5752 ( .A(datapointV_1_fu_674_p2[4]), .B(n397), .Y(n411) );
  INVX1 U5753 ( .A(n411), .Y(n5193) );
  AND2X1 U5754 ( .A(datapointV_1_fu_674_p2[5]), .B(n397), .Y(n409) );
  INVX1 U5755 ( .A(n409), .Y(n5194) );
  AND2X1 U5756 ( .A(datapointV_1_fu_674_p2[6]), .B(n397), .Y(n407) );
  INVX1 U5757 ( .A(n407), .Y(n5195) );
  AND2X1 U5758 ( .A(datapointV_1_fu_674_p2[7]), .B(n397), .Y(n405) );
  INVX1 U5759 ( .A(n405), .Y(n5196) );
  AND2X1 U5760 ( .A(datapointV_1_fu_674_p2[8]), .B(n397), .Y(n403) );
  INVX1 U5761 ( .A(n403), .Y(n5197) );
  AND2X1 U5762 ( .A(datapointV_1_fu_674_p2[9]), .B(n397), .Y(n401) );
  INVX1 U5763 ( .A(n401), .Y(n5198) );
  BUFX2 U5764 ( .A(\Decision_AXILiteS_s_axi_U/n646 ), .Y(n5199) );
  AND2X1 U5765 ( .A(\recentABools_data_q0[0] ), .B(N461), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n17 ) );
  INVX1 U5766 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n17 ), 
        .Y(n5200) );
  AND2X1 U5767 ( .A(\recentVBools_data_q0[0] ), .B(N466), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n16 ) );
  INVX1 U5768 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n16 ), 
        .Y(n5201) );
  AND2X1 U5769 ( .A(ACaptureThresh_loc_reg_288[0]), .B(n8969), .Y(n3062) );
  INVX1 U5770 ( .A(n3062), .Y(n5202) );
  AND2X1 U5771 ( .A(ACaptureThresh_loc_reg_288[1]), .B(n8970), .Y(n3060) );
  INVX1 U5772 ( .A(n3060), .Y(n5203) );
  AND2X1 U5773 ( .A(ACaptureThresh_loc_reg_288[2]), .B(n8971), .Y(n3058) );
  INVX1 U5774 ( .A(n3058), .Y(n5204) );
  BUFX2 U5775 ( .A(n3061), .Y(n5205) );
  BUFX2 U5776 ( .A(n3059), .Y(n5206) );
  BUFX2 U5777 ( .A(n3057), .Y(n5207) );
  BUFX2 U5778 ( .A(n11168), .Y(n5208) );
  BUFX2 U5779 ( .A(n11545), .Y(n5209) );
  BUFX2 U5780 ( .A(n11714), .Y(n5210) );
  BUFX2 U5781 ( .A(n11803), .Y(n5211) );
  BUFX2 U5782 ( .A(n11892), .Y(n5212) );
  BUFX2 U5783 ( .A(n12000), .Y(n5213) );
  BUFX2 U5784 ( .A(n12089), .Y(n5214) );
  BUFX2 U5785 ( .A(n12178), .Y(n5215) );
  BUFX2 U5786 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n16 ), 
        .Y(n5216) );
  BUFX2 U5787 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n15 ), 
        .Y(n5217) );
  BUFX2 U5788 ( .A(\Decision_AXILiteS_s_axi_U/n626 ), .Y(n5218) );
  BUFX2 U5789 ( .A(\Decision_AXILiteS_s_axi_U/n645 ), .Y(n5219) );
  AND2X1 U5790 ( .A(s_axi_AXILiteS_RDATA[7]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n249 ) );
  INVX1 U5791 ( .A(\Decision_AXILiteS_s_axi_U/n249 ), .Y(n5220) );
  AND2X1 U5792 ( .A(s_axi_AXILiteS_RDATA[3]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n279 ) );
  INVX1 U5793 ( .A(\Decision_AXILiteS_s_axi_U/n279 ), .Y(n5221) );
  AND2X1 U5794 ( .A(s_axi_AXILiteS_RDATA[2]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n288 ) );
  INVX1 U5795 ( .A(\Decision_AXILiteS_s_axi_U/n288 ), .Y(n5222) );
  AND2X1 U5796 ( .A(s_axi_AXILiteS_RDATA[1]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n297 ) );
  INVX1 U5797 ( .A(\Decision_AXILiteS_s_axi_U/n297 ), .Y(n5223) );
  AND2X1 U5798 ( .A(s_axi_AXILiteS_RDATA[0]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n311 ) );
  INVX1 U5799 ( .A(\Decision_AXILiteS_s_axi_U/n311 ), .Y(n5224) );
  BUFX2 U5800 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n9 ), 
        .Y(n5225) );
  BUFX2 U5801 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n14 ), 
        .Y(n5226) );
  BUFX2 U5802 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n8 ), 
        .Y(n5227) );
  BUFX2 U5803 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n26 ), 
        .Y(n5228) );
  BUFX2 U5804 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n50 ), 
        .Y(n5229) );
  BUFX2 U5805 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n58 ), 
        .Y(n5230) );
  BUFX2 U5806 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n71 ), 
        .Y(n5231) );
  BUFX2 U5807 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n79 ), 
        .Y(n5232) );
  BUFX2 U5808 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n92 ), 
        .Y(n5233) );
  BUFX2 U5809 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n100 ), 
        .Y(n5234) );
  BUFX2 U5810 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n113 ), 
        .Y(n5235) );
  BUFX2 U5811 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n121 ), 
        .Y(n5236) );
  BUFX2 U5812 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n134 ), 
        .Y(n5237) );
  BUFX2 U5813 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n142 ), 
        .Y(n5238) );
  BUFX2 U5814 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n155 ), 
        .Y(n5239) );
  BUFX2 U5815 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n163 ), 
        .Y(n5240) );
  BUFX2 U5816 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n176 ), 
        .Y(n5241) );
  BUFX2 U5817 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n184 ), 
        .Y(n5242) );
  BUFX2 U5818 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n197 ), 
        .Y(n5243) );
  BUFX2 U5819 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n205 ), 
        .Y(n5244) );
  BUFX2 U5820 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n218 ), 
        .Y(n5245) );
  BUFX2 U5821 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n226 ), 
        .Y(n5246) );
  BUFX2 U5822 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n239 ), 
        .Y(n5247) );
  BUFX2 U5823 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n247 ), 
        .Y(n5248) );
  BUFX2 U5824 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n260 ), 
        .Y(n5249) );
  BUFX2 U5825 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n268 ), 
        .Y(n5250) );
  BUFX2 U5826 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n281 ), 
        .Y(n5251) );
  BUFX2 U5827 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n289 ), 
        .Y(n5252) );
  BUFX2 U5828 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n302 ), 
        .Y(n5253) );
  BUFX2 U5829 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n310 ), 
        .Y(n5254) );
  BUFX2 U5830 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n323 ), 
        .Y(n5255) );
  BUFX2 U5831 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n331 ), 
        .Y(n5256) );
  BUFX2 U5832 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n344 ), 
        .Y(n5257) );
  BUFX2 U5833 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n355 ), 
        .Y(n5258) );
  BUFX2 U5834 ( .A(n1932), .Y(n5259) );
  BUFX2 U5835 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n9 ), 
        .Y(n5260) );
  BUFX2 U5836 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n27 ), 
        .Y(n5261) );
  BUFX2 U5837 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n51 ), 
        .Y(n5262) );
  BUFX2 U5838 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n59 ), 
        .Y(n5263) );
  BUFX2 U5839 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n72 ), 
        .Y(n5264) );
  BUFX2 U5840 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n80 ), 
        .Y(n5265) );
  BUFX2 U5841 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n93 ), 
        .Y(n5266) );
  BUFX2 U5842 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n101 ), 
        .Y(n5267) );
  BUFX2 U5843 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n114 ), 
        .Y(n5268) );
  BUFX2 U5844 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n122 ), 
        .Y(n5269) );
  BUFX2 U5845 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n135 ), 
        .Y(n5270) );
  BUFX2 U5846 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n143 ), 
        .Y(n5271) );
  BUFX2 U5847 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n156 ), 
        .Y(n5272) );
  BUFX2 U5848 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n164 ), 
        .Y(n5273) );
  BUFX2 U5849 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n177 ), 
        .Y(n5274) );
  BUFX2 U5850 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n185 ), 
        .Y(n5275) );
  BUFX2 U5851 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n198 ), 
        .Y(n5276) );
  BUFX2 U5852 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n206 ), 
        .Y(n5277) );
  BUFX2 U5853 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n219 ), 
        .Y(n5278) );
  BUFX2 U5854 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n227 ), 
        .Y(n5279) );
  BUFX2 U5855 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n240 ), 
        .Y(n5280) );
  BUFX2 U5856 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n248 ), 
        .Y(n5281) );
  BUFX2 U5857 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n261 ), 
        .Y(n5282) );
  BUFX2 U5858 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n269 ), 
        .Y(n5283) );
  BUFX2 U5859 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n282 ), 
        .Y(n5284) );
  BUFX2 U5860 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n290 ), 
        .Y(n5285) );
  BUFX2 U5861 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n303 ), 
        .Y(n5286) );
  BUFX2 U5862 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n311 ), 
        .Y(n5287) );
  BUFX2 U5863 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n324 ), 
        .Y(n5288) );
  BUFX2 U5864 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n332 ), 
        .Y(n5289) );
  BUFX2 U5865 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n345 ), 
        .Y(n5290) );
  BUFX2 U5866 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n356 ), 
        .Y(n5291) );
  BUFX2 U5867 ( .A(n1933), .Y(n5292) );
  BUFX2 U5868 ( .A(\Decision_AXILiteS_s_axi_U/n459 ), .Y(n5293) );
  BUFX2 U5869 ( .A(\Decision_AXILiteS_s_axi_U/n566 ), .Y(n5294) );
  BUFX2 U5870 ( .A(n11122), .Y(n5295) );
  BUFX2 U5871 ( .A(n11499), .Y(n5296) );
  BUFX2 U5872 ( .A(n11543), .Y(n5297) );
  BUFX2 U5873 ( .A(n11668), .Y(n5298) );
  BUFX2 U5874 ( .A(n11712), .Y(n5299) );
  BUFX2 U5875 ( .A(n11757), .Y(n5300) );
  BUFX2 U5876 ( .A(n11801), .Y(n5301) );
  BUFX2 U5877 ( .A(n11846), .Y(n5302) );
  BUFX2 U5878 ( .A(n11954), .Y(n5303) );
  BUFX2 U5879 ( .A(n11998), .Y(n5304) );
  BUFX2 U5880 ( .A(n12043), .Y(n5305) );
  BUFX2 U5881 ( .A(n12087), .Y(n5306) );
  BUFX2 U5882 ( .A(n12132), .Y(n5307) );
  BUFX2 U5883 ( .A(n12176), .Y(n5308) );
  BUFX2 U5884 ( .A(n11261), .Y(n5309) );
  BUFX2 U5885 ( .A(n11265), .Y(n5310) );
  BUFX2 U5886 ( .A(n11269), .Y(n5311) );
  BUFX2 U5887 ( .A(n11273), .Y(n5312) );
  BUFX2 U5888 ( .A(n11277), .Y(n5313) );
  BUFX2 U5889 ( .A(n11281), .Y(n5314) );
  BUFX2 U5890 ( .A(n11285), .Y(n5315) );
  BUFX2 U5891 ( .A(n11289), .Y(n5316) );
  BUFX2 U5892 ( .A(n11293), .Y(n5317) );
  BUFX2 U5893 ( .A(n11297), .Y(n5318) );
  BUFX2 U5894 ( .A(n11301), .Y(n5319) );
  BUFX2 U5895 ( .A(n11313), .Y(n5320) );
  BUFX2 U5896 ( .A(n11317), .Y(n5321) );
  BUFX2 U5897 ( .A(n11321), .Y(n5322) );
  BUFX2 U5898 ( .A(n11325), .Y(n5323) );
  BUFX2 U5899 ( .A(n11329), .Y(n5324) );
  BUFX2 U5900 ( .A(n11333), .Y(n5325) );
  BUFX2 U5901 ( .A(n11337), .Y(n5326) );
  BUFX2 U5902 ( .A(n11341), .Y(n5327) );
  BUFX2 U5903 ( .A(n11345), .Y(n5328) );
  BUFX2 U5904 ( .A(n11349), .Y(n5329) );
  BUFX2 U5905 ( .A(n11353), .Y(n5330) );
  BUFX2 U5906 ( .A(n11365), .Y(n5331) );
  BUFX2 U5907 ( .A(n11369), .Y(n5332) );
  BUFX2 U5908 ( .A(n11373), .Y(n5333) );
  BUFX2 U5909 ( .A(n11377), .Y(n5334) );
  BUFX2 U5910 ( .A(n11381), .Y(n5335) );
  BUFX2 U5911 ( .A(n11385), .Y(n5336) );
  BUFX2 U5912 ( .A(n11389), .Y(n5337) );
  BUFX2 U5913 ( .A(n11393), .Y(n5338) );
  BUFX2 U5914 ( .A(n11397), .Y(n5339) );
  BUFX2 U5915 ( .A(n11401), .Y(n5340) );
  BUFX2 U5916 ( .A(n11405), .Y(n5341) );
  BUFX2 U5917 ( .A(n11417), .Y(n5342) );
  BUFX2 U5918 ( .A(n11421), .Y(n5343) );
  BUFX2 U5919 ( .A(n11425), .Y(n5344) );
  BUFX2 U5920 ( .A(n11429), .Y(n5345) );
  BUFX2 U5921 ( .A(n11433), .Y(n5346) );
  BUFX2 U5922 ( .A(n11437), .Y(n5347) );
  BUFX2 U5923 ( .A(n11441), .Y(n5348) );
  BUFX2 U5924 ( .A(n11445), .Y(n5349) );
  BUFX2 U5925 ( .A(n11449), .Y(n5350) );
  BUFX2 U5926 ( .A(n11453), .Y(n5351) );
  BUFX2 U5927 ( .A(n11457), .Y(n5352) );
  BUFX2 U5928 ( .A(n11612), .Y(n5353) );
  BUFX2 U5929 ( .A(n12245), .Y(n5354) );
  BUFX2 U5930 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n10 ), 
        .Y(n5355) );
  BUFX2 U5931 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n18 ), 
        .Y(n5356) );
  BUFX2 U5932 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n28 ), 
        .Y(n5357) );
  BUFX2 U5933 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n36 ), 
        .Y(n5358) );
  BUFX2 U5934 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n52 ), 
        .Y(n5359) );
  BUFX2 U5935 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n55 ), 
        .Y(n5360) );
  BUFX2 U5936 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n60 ), 
        .Y(n5361) );
  BUFX2 U5937 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n63 ), 
        .Y(n5362) );
  BUFX2 U5938 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n73 ), 
        .Y(n5363) );
  BUFX2 U5939 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n76 ), 
        .Y(n5364) );
  BUFX2 U5940 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n81 ), 
        .Y(n5365) );
  BUFX2 U5941 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n84 ), 
        .Y(n5366) );
  BUFX2 U5942 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n94 ), 
        .Y(n5367) );
  BUFX2 U5943 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n97 ), 
        .Y(n5368) );
  BUFX2 U5944 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n102 ), 
        .Y(n5369) );
  BUFX2 U5945 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n105 ), 
        .Y(n5370) );
  BUFX2 U5946 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n115 ), 
        .Y(n5371) );
  BUFX2 U5947 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n118 ), 
        .Y(n5372) );
  BUFX2 U5948 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n123 ), 
        .Y(n5373) );
  BUFX2 U5949 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n126 ), 
        .Y(n5374) );
  BUFX2 U5950 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n136 ), 
        .Y(n5375) );
  BUFX2 U5951 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n139 ), 
        .Y(n5376) );
  BUFX2 U5952 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n144 ), 
        .Y(n5377) );
  BUFX2 U5953 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n147 ), 
        .Y(n5378) );
  BUFX2 U5954 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n157 ), 
        .Y(n5379) );
  BUFX2 U5955 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n160 ), 
        .Y(n5380) );
  BUFX2 U5956 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n165 ), 
        .Y(n5381) );
  BUFX2 U5957 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n168 ), 
        .Y(n5382) );
  BUFX2 U5958 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n178 ), 
        .Y(n5383) );
  BUFX2 U5959 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n181 ), 
        .Y(n5384) );
  BUFX2 U5960 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n186 ), 
        .Y(n5385) );
  BUFX2 U5961 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n189 ), 
        .Y(n5386) );
  BUFX2 U5962 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n199 ), 
        .Y(n5387) );
  BUFX2 U5963 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n202 ), 
        .Y(n5388) );
  BUFX2 U5964 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n207 ), 
        .Y(n5389) );
  BUFX2 U5965 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n210 ), 
        .Y(n5390) );
  BUFX2 U5966 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n220 ), 
        .Y(n5391) );
  BUFX2 U5967 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n223 ), 
        .Y(n5392) );
  BUFX2 U5968 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n228 ), 
        .Y(n5393) );
  BUFX2 U5969 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n231 ), 
        .Y(n5394) );
  BUFX2 U5970 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n241 ), 
        .Y(n5395) );
  BUFX2 U5971 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n244 ), 
        .Y(n5396) );
  BUFX2 U5972 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n249 ), 
        .Y(n5397) );
  BUFX2 U5973 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n252 ), 
        .Y(n5398) );
  BUFX2 U5974 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n262 ), 
        .Y(n5399) );
  BUFX2 U5975 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n265 ), 
        .Y(n5400) );
  BUFX2 U5976 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n270 ), 
        .Y(n5401) );
  BUFX2 U5977 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n273 ), 
        .Y(n5402) );
  BUFX2 U5978 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n283 ), 
        .Y(n5403) );
  BUFX2 U5979 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n286 ), 
        .Y(n5404) );
  BUFX2 U5980 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n291 ), 
        .Y(n5405) );
  BUFX2 U5981 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n294 ), 
        .Y(n5406) );
  BUFX2 U5982 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n304 ), 
        .Y(n5407) );
  BUFX2 U5983 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n307 ), 
        .Y(n5408) );
  BUFX2 U5984 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n312 ), 
        .Y(n5409) );
  BUFX2 U5985 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n315 ), 
        .Y(n5410) );
  BUFX2 U5986 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n325 ), 
        .Y(n5411) );
  BUFX2 U5987 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n328 ), 
        .Y(n5412) );
  BUFX2 U5988 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n333 ), 
        .Y(n5413) );
  BUFX2 U5989 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n336 ), 
        .Y(n5414) );
  BUFX2 U5990 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n346 ), 
        .Y(n5415) );
  BUFX2 U5991 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n349 ), 
        .Y(n5416) );
  BUFX2 U5992 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n357 ), 
        .Y(n5417) );
  BUFX2 U5993 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n367 ), 
        .Y(n5418) );
  BUFX2 U5994 ( .A(\Decision_AXILiteS_s_axi_U/n152 ), .Y(n5419) );
  BUFX2 U5995 ( .A(\Decision_AXILiteS_s_axi_U/n160 ), .Y(n5420) );
  BUFX2 U5996 ( .A(\Decision_AXILiteS_s_axi_U/n163 ), .Y(n5421) );
  BUFX2 U5997 ( .A(\Decision_AXILiteS_s_axi_U/n166 ), .Y(n5422) );
  BUFX2 U5998 ( .A(\Decision_AXILiteS_s_axi_U/n169 ), .Y(n5423) );
  BUFX2 U5999 ( .A(\Decision_AXILiteS_s_axi_U/n172 ), .Y(n5424) );
  BUFX2 U6000 ( .A(\Decision_AXILiteS_s_axi_U/n175 ), .Y(n5425) );
  BUFX2 U6001 ( .A(\Decision_AXILiteS_s_axi_U/n178 ), .Y(n5426) );
  BUFX2 U6002 ( .A(\Decision_AXILiteS_s_axi_U/n181 ), .Y(n5427) );
  BUFX2 U6003 ( .A(\Decision_AXILiteS_s_axi_U/n184 ), .Y(n5428) );
  BUFX2 U6004 ( .A(\Decision_AXILiteS_s_axi_U/n187 ), .Y(n5429) );
  BUFX2 U6005 ( .A(\Decision_AXILiteS_s_axi_U/n190 ), .Y(n5430) );
  BUFX2 U6006 ( .A(\Decision_AXILiteS_s_axi_U/n193 ), .Y(n5431) );
  BUFX2 U6007 ( .A(\Decision_AXILiteS_s_axi_U/n196 ), .Y(n5432) );
  BUFX2 U6008 ( .A(\Decision_AXILiteS_s_axi_U/n199 ), .Y(n5433) );
  BUFX2 U6009 ( .A(\Decision_AXILiteS_s_axi_U/n202 ), .Y(n5434) );
  BUFX2 U6010 ( .A(\Decision_AXILiteS_s_axi_U/n205 ), .Y(n5435) );
  BUFX2 U6011 ( .A(\Decision_AXILiteS_s_axi_U/n212 ), .Y(n5436) );
  BUFX2 U6012 ( .A(\Decision_AXILiteS_s_axi_U/n217 ), .Y(n5437) );
  BUFX2 U6013 ( .A(\Decision_AXILiteS_s_axi_U/n222 ), .Y(n5438) );
  BUFX2 U6014 ( .A(\Decision_AXILiteS_s_axi_U/n227 ), .Y(n5439) );
  BUFX2 U6015 ( .A(\Decision_AXILiteS_s_axi_U/n232 ), .Y(n5440) );
  BUFX2 U6016 ( .A(\Decision_AXILiteS_s_axi_U/n237 ), .Y(n5441) );
  BUFX2 U6017 ( .A(\Decision_AXILiteS_s_axi_U/n242 ), .Y(n5442) );
  BUFX2 U6018 ( .A(\Decision_AXILiteS_s_axi_U/n255 ), .Y(n5443) );
  BUFX2 U6019 ( .A(\Decision_AXILiteS_s_axi_U/n260 ), .Y(n5444) );
  BUFX2 U6020 ( .A(\Decision_AXILiteS_s_axi_U/n267 ), .Y(n5445) );
  BUFX2 U6021 ( .A(\Decision_AXILiteS_s_axi_U/n274 ), .Y(n5446) );
  BUFX2 U6022 ( .A(\Decision_AXILiteS_s_axi_U/n285 ), .Y(n5447) );
  BUFX2 U6023 ( .A(\Decision_AXILiteS_s_axi_U/n294 ), .Y(n5448) );
  BUFX2 U6024 ( .A(\Decision_AXILiteS_s_axi_U/n326 ), .Y(n5449) );
  BUFX2 U6025 ( .A(n361), .Y(n5450) );
  BUFX2 U6026 ( .A(n358), .Y(n5451) );
  BUFX2 U6027 ( .A(n11099), .Y(n5452) );
  BUFX2 U6028 ( .A(n11139), .Y(n5453) );
  BUFX2 U6029 ( .A(n11146), .Y(n5454) );
  BUFX2 U6030 ( .A(n11476), .Y(n5455) );
  BUFX2 U6031 ( .A(n11516), .Y(n5456) );
  BUFX2 U6032 ( .A(n11524), .Y(n5457) );
  BUFX2 U6033 ( .A(n11601), .Y(n5458) );
  BUFX2 U6034 ( .A(n11578), .Y(n5459) );
  BUFX2 U6035 ( .A(n11594), .Y(n5460) );
  BUFX2 U6036 ( .A(n11645), .Y(n5461) );
  BUFX2 U6037 ( .A(n11685), .Y(n5462) );
  BUFX2 U6038 ( .A(n11692), .Y(n5463) );
  BUFX2 U6039 ( .A(n11734), .Y(n5464) );
  BUFX2 U6040 ( .A(n11774), .Y(n5465) );
  BUFX2 U6041 ( .A(n11782), .Y(n5466) );
  BUFX2 U6042 ( .A(n11823), .Y(n5467) );
  BUFX2 U6043 ( .A(n11863), .Y(n5468) );
  BUFX2 U6044 ( .A(n11870), .Y(n5469) );
  BUFX2 U6045 ( .A(n11931), .Y(n5470) );
  BUFX2 U6046 ( .A(n11971), .Y(n5471) );
  BUFX2 U6047 ( .A(n11978), .Y(n5472) );
  BUFX2 U6048 ( .A(n12020), .Y(n5473) );
  BUFX2 U6049 ( .A(n12060), .Y(n5474) );
  BUFX2 U6050 ( .A(n12067), .Y(n5475) );
  BUFX2 U6051 ( .A(n12109), .Y(n5476) );
  BUFX2 U6052 ( .A(n12149), .Y(n5477) );
  BUFX2 U6053 ( .A(n12156), .Y(n5478) );
  BUFX2 U6054 ( .A(n12234), .Y(n5479) );
  BUFX2 U6055 ( .A(n12211), .Y(n5480) );
  BUFX2 U6056 ( .A(n12227), .Y(n5481) );
  BUFX2 U6057 ( .A(\Decision_AXILiteS_s_axi_U/n304 ), .Y(n5482) );
  BUFX2 U6058 ( .A(\Decision_AXILiteS_s_axi_U/n595 ), .Y(n5483) );
  AND2X1 U6059 ( .A(data_read_reg_1495[0]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1 )
         );
  INVX1 U6060 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n1 ), 
        .Y(n5484) );
  AND2X1 U6061 ( .A(data_read_reg_1495[1]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n45 )
         );
  INVX1 U6062 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n45 ), 
        .Y(n5485) );
  AND2X1 U6063 ( .A(data_read_reg_1495[2]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n66 )
         );
  INVX1 U6064 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n66 ), 
        .Y(n5486) );
  AND2X1 U6065 ( .A(data_read_reg_1495[3]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n87 )
         );
  INVX1 U6066 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n87 ), 
        .Y(n5487) );
  AND2X1 U6067 ( .A(data_read_reg_1495[4]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n108 ) );
  INVX1 U6068 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n108 ), 
        .Y(n5488) );
  AND2X1 U6069 ( .A(data_read_reg_1495[5]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n129 ) );
  INVX1 U6070 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n129 ), 
        .Y(n5489) );
  AND2X1 U6071 ( .A(data_read_reg_1495[6]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n150 ) );
  INVX1 U6072 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n150 ), 
        .Y(n5490) );
  AND2X1 U6073 ( .A(data_read_reg_1495[7]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n171 ) );
  INVX1 U6074 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n171 ), 
        .Y(n5491) );
  AND2X1 U6075 ( .A(data_read_reg_1495[8]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n192 ) );
  INVX1 U6076 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n192 ), 
        .Y(n5492) );
  AND2X1 U6077 ( .A(data_read_reg_1495[9]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n213 ) );
  INVX1 U6078 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n213 ), 
        .Y(n5493) );
  AND2X1 U6079 ( .A(data_read_reg_1495[10]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n234 ) );
  INVX1 U6080 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n234 ), 
        .Y(n5494) );
  AND2X1 U6081 ( .A(data_read_reg_1495[11]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n255 ) );
  INVX1 U6082 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n255 ), 
        .Y(n5495) );
  AND2X1 U6083 ( .A(data_read_reg_1495[12]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n276 ) );
  INVX1 U6084 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n276 ), 
        .Y(n5496) );
  AND2X1 U6085 ( .A(data_read_reg_1495[13]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n297 ) );
  INVX1 U6086 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n297 ), 
        .Y(n5497) );
  AND2X1 U6087 ( .A(data_read_reg_1495[14]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n318 ) );
  INVX1 U6088 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n318 ), 
        .Y(n5498) );
  AND2X1 U6089 ( .A(data_read_reg_1495[15]), .B(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n339 ) );
  INVX1 U6090 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n339 ), 
        .Y(n5499) );
  AND2X1 U6091 ( .A(ap_rst_n), .B(ap_CS_fsm[13]), .Y(
        \Decision_AXILiteS_s_axi_U/n620 ) );
  INVX1 U6092 ( .A(\Decision_AXILiteS_s_axi_U/n620 ), .Y(n5500) );
  BUFX2 U6093 ( .A(n11123), .Y(n5501) );
  BUFX2 U6094 ( .A(n11500), .Y(n5502) );
  BUFX2 U6095 ( .A(n11607), .Y(n5503) );
  BUFX2 U6096 ( .A(n11669), .Y(n5504) );
  BUFX2 U6097 ( .A(n11758), .Y(n5505) );
  BUFX2 U6098 ( .A(n11847), .Y(n5506) );
  BUFX2 U6099 ( .A(n11955), .Y(n5507) );
  BUFX2 U6100 ( .A(n12044), .Y(n5508) );
  BUFX2 U6101 ( .A(n12133), .Y(n5509) );
  BUFX2 U6102 ( .A(n12240), .Y(n5510) );
  BUFX2 U6103 ( .A(n11488), .Y(n5511) );
  BUFX2 U6104 ( .A(n11544), .Y(n5512) );
  BUFX2 U6105 ( .A(n11657), .Y(n5513) );
  BUFX2 U6106 ( .A(n11713), .Y(n5514) );
  BUFX2 U6107 ( .A(n11746), .Y(n5515) );
  BUFX2 U6108 ( .A(n11802), .Y(n5516) );
  BUFX2 U6109 ( .A(n11943), .Y(n5517) );
  BUFX2 U6110 ( .A(n11999), .Y(n5518) );
  BUFX2 U6111 ( .A(n12121), .Y(n5519) );
  BUFX2 U6112 ( .A(n12177), .Y(n5520) );
  BUFX2 U6113 ( .A(n11076), .Y(n5521) );
  BUFX2 U6114 ( .A(n11124), .Y(n5522) );
  BUFX2 U6115 ( .A(n11501), .Y(n5523) );
  BUFX2 U6116 ( .A(n11670), .Y(n5524) );
  BUFX2 U6117 ( .A(n11759), .Y(n5525) );
  BUFX2 U6118 ( .A(n11848), .Y(n5526) );
  BUFX2 U6119 ( .A(n11956), .Y(n5527) );
  BUFX2 U6120 ( .A(n12045), .Y(n5528) );
  BUFX2 U6121 ( .A(n12134), .Y(n5529) );
  BUFX2 U6122 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n1 ), 
        .Y(n5530) );
  BUFX2 U6123 ( .A(\Decision_AXILiteS_s_axi_U/n336 ), .Y(n5531) );
  BUFX2 U6124 ( .A(\Decision_AXILiteS_s_axi_U/n618 ), .Y(n5532) );
  BUFX2 U6125 ( .A(n11174), .Y(n5533) );
  BUFX2 U6126 ( .A(n11551), .Y(n5534) );
  BUFX2 U6127 ( .A(n11628), .Y(n5535) );
  BUFX2 U6128 ( .A(n11720), .Y(n5536) );
  BUFX2 U6129 ( .A(n11809), .Y(n5537) );
  BUFX2 U6130 ( .A(n11898), .Y(n5538) );
  BUFX2 U6131 ( .A(n12006), .Y(n5539) );
  BUFX2 U6132 ( .A(n12095), .Y(n5540) );
  BUFX2 U6133 ( .A(n12184), .Y(n5541) );
  BUFX2 U6134 ( .A(n12261), .Y(n5542) );
  BUFX2 U6135 ( .A(\Decision_AXILiteS_s_axi_U/n251 ), .Y(n5543) );
  BUFX2 U6136 ( .A(\Decision_AXILiteS_s_axi_U/n281 ), .Y(n5544) );
  BUFX2 U6137 ( .A(\Decision_AXILiteS_s_axi_U/n290 ), .Y(n5545) );
  BUFX2 U6138 ( .A(\Decision_AXILiteS_s_axi_U/n299 ), .Y(n5546) );
  BUFX2 U6139 ( .A(\Decision_AXILiteS_s_axi_U/n313 ), .Y(n5547) );
  BUFX2 U6140 ( .A(n1649), .Y(n5548) );
  AND2X1 U6141 ( .A(n7779), .B(n7569), .Y(n11631) );
  INVX1 U6142 ( .A(n11631), .Y(n5549) );
  AND2X1 U6143 ( .A(n7777), .B(n7567), .Y(n12264) );
  INVX1 U6144 ( .A(n12264), .Y(n5550) );
  BUFX2 U6145 ( .A(n11126), .Y(n5551) );
  BUFX2 U6146 ( .A(n11503), .Y(n5552) );
  BUFX2 U6147 ( .A(n11672), .Y(n5553) );
  BUFX2 U6148 ( .A(n11761), .Y(n5554) );
  BUFX2 U6149 ( .A(n11850), .Y(n5555) );
  BUFX2 U6150 ( .A(n11958), .Y(n5556) );
  BUFX2 U6151 ( .A(n12047), .Y(n5557) );
  BUFX2 U6152 ( .A(n12136), .Y(n5558) );
  BUFX2 U6153 ( .A(\Decision_AXILiteS_s_axi_U/n259 ), .Y(n5559) );
  BUFX2 U6154 ( .A(\Decision_AXILiteS_s_axi_U/n266 ), .Y(n5560) );
  BUFX2 U6155 ( .A(\Decision_AXILiteS_s_axi_U/n273 ), .Y(n5561) );
  BUFX2 U6156 ( .A(n11066), .Y(n5562) );
  BUFX2 U6157 ( .A(n11084), .Y(n5563) );
  BUFX2 U6158 ( .A(\Decision_AXILiteS_s_axi_U/n261 ), .Y(n5564) );
  BUFX2 U6159 ( .A(\Decision_AXILiteS_s_axi_U/n268 ), .Y(n5565) );
  BUFX2 U6160 ( .A(\Decision_AXILiteS_s_axi_U/n275 ), .Y(n5566) );
  BUFX2 U6161 ( .A(n11609), .Y(n5567) );
  BUFX2 U6162 ( .A(n12242), .Y(n5568) );
  BUFX2 U6163 ( .A(\Decision_AXILiteS_s_axi_U/n596 ), .Y(n5569) );
  BUFX2 U6164 ( .A(\Decision_AXILiteS_s_axi_U/n628 ), .Y(n5570) );
  AND2X1 U6165 ( .A(VbeatDelay_new_1_reg_326[25]), .B(n10729), .Y(n11138) );
  INVX1 U6166 ( .A(n11138), .Y(n5571) );
  AND2X1 U6167 ( .A(sum_phi_fu_311_p4[9]), .B(n9683), .Y(n11469) );
  INVX1 U6168 ( .A(n11469), .Y(n5572) );
  AND2X1 U6169 ( .A(sum_phi_fu_311_p4[13]), .B(n9699), .Y(n11475) );
  INVX1 U6170 ( .A(n11475), .Y(n5573) );
  AND2X1 U6171 ( .A(sum_phi_fu_311_p4[25]), .B(n9747), .Y(n11515) );
  INVX1 U6172 ( .A(n11515), .Y(n5574) );
  AND2X1 U6173 ( .A(sum_phi_fu_311_p4[29]), .B(n9761), .Y(n11523) );
  INVX1 U6174 ( .A(n11523), .Y(n5575) );
  INVX1 U6175 ( .A(n11573), .Y(n5576) );
  AND2X1 U6176 ( .A(p_1_cast_fu_1031_p1[5]), .B(n9769), .Y(n11577) );
  INVX1 U6177 ( .A(n11577), .Y(n5577) );
  AND2X1 U6178 ( .A(p_1_cast_fu_1031_p1[9]), .B(n9771), .Y(n11587) );
  INVX1 U6179 ( .A(n11587), .Y(n5578) );
  AND2X1 U6180 ( .A(p_1_cast_fu_1031_p1[13]), .B(n9774), .Y(n11593) );
  INVX1 U6181 ( .A(n11593), .Y(n5579) );
  AND2X1 U6182 ( .A(p_1_cast_fu_1031_p1_31), .B(n9779), .Y(n11611) );
  INVX1 U6183 ( .A(n11611), .Y(n5580) );
  AND2X1 U6184 ( .A(p_1_cast_fu_1031_p1_31), .B(n9782), .Y(n11625) );
  INVX1 U6185 ( .A(n11625), .Y(n5581) );
  AND2X1 U6186 ( .A(n2275), .B(n9586), .Y(n11644) );
  INVX1 U6187 ( .A(n11644), .Y(n5582) );
  AND2X1 U6188 ( .A(n2251), .B(n9626), .Y(n11684) );
  INVX1 U6189 ( .A(n11684), .Y(n5583) );
  AND2X1 U6190 ( .A(n2243), .B(n9638), .Y(n11691) );
  INVX1 U6191 ( .A(n11691), .Y(n5584) );
  AND2X1 U6192 ( .A(sum_1_phi_fu_379_p4[9]), .B(n9579), .Y(n11727) );
  INVX1 U6193 ( .A(n11727), .Y(n5585) );
  AND2X1 U6194 ( .A(sum_1_phi_fu_379_p4[13]), .B(n9592), .Y(n11733) );
  INVX1 U6195 ( .A(n11733), .Y(n5586) );
  AND2X1 U6196 ( .A(sum_1_phi_fu_379_p4[25]), .B(n9632), .Y(n11773) );
  INVX1 U6197 ( .A(n11773), .Y(n5587) );
  AND2X1 U6198 ( .A(sum_1_phi_fu_379_p4[29]), .B(n9644), .Y(n11781) );
  INVX1 U6199 ( .A(n11781), .Y(n5588) );
  AND2X1 U6200 ( .A(VbeatDelay_new_1_reg_326[25]), .B(n10433), .Y(n11862) );
  INVX1 U6201 ( .A(n11862), .Y(n5589) );
  AND2X1 U6202 ( .A(tmp_6_reg_1538[25]), .B(n9626), .Y(n11970) );
  INVX1 U6203 ( .A(n11970), .Y(n5590) );
  AND2X1 U6204 ( .A(tmp_7_reg_1544[25]), .B(n9741), .Y(n12059) );
  INVX1 U6205 ( .A(n12059), .Y(n5591) );
  AND2X1 U6206 ( .A(n2768), .B(n9693), .Y(n12108) );
  INVX1 U6207 ( .A(n12108), .Y(n5592) );
  AND2X1 U6208 ( .A(n2744), .B(n9741), .Y(n12148) );
  INVX1 U6209 ( .A(n12148), .Y(n5593) );
  AND2X1 U6210 ( .A(n2736), .B(n9755), .Y(n12155) );
  INVX1 U6211 ( .A(n12155), .Y(n5594) );
  INVX1 U6212 ( .A(n12206), .Y(n5595) );
  AND2X1 U6213 ( .A(p_cast_fu_688_p1[5]), .B(n9501), .Y(n12210) );
  INVX1 U6214 ( .A(n12210), .Y(n5596) );
  AND2X1 U6215 ( .A(p_cast_fu_688_p1[9]), .B(n9507), .Y(n12220) );
  INVX1 U6216 ( .A(n12220), .Y(n5597) );
  AND2X1 U6217 ( .A(p_cast_fu_688_p1[13]), .B(n9513), .Y(n12226) );
  INVX1 U6218 ( .A(n12226), .Y(n5598) );
  AND2X1 U6219 ( .A(p_cast_fu_688_p1_31), .B(n9520), .Y(n12244) );
  INVX1 U6220 ( .A(n12244), .Y(n5599) );
  AND2X1 U6221 ( .A(p_cast_fu_688_p1_31), .B(n9523), .Y(n12258) );
  INVX1 U6222 ( .A(n12258), .Y(n5600) );
  AND2X1 U6223 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][0] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n11 ) );
  INVX1 U6224 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n11 ), 
        .Y(n5601) );
  AND2X1 U6225 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][0] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n19 ) );
  INVX1 U6226 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n19 ), 
        .Y(n5602) );
  AND2X1 U6227 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][0] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n29 ) );
  INVX1 U6228 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n29 ), 
        .Y(n5603) );
  AND2X1 U6229 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][0] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n37 ) );
  INVX1 U6230 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n37 ), 
        .Y(n5604) );
  AND2X1 U6231 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][1] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n53 ) );
  INVX1 U6232 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n53 ), 
        .Y(n5605) );
  AND2X1 U6233 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][1] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n56 ) );
  INVX1 U6234 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n56 ), 
        .Y(n5606) );
  AND2X1 U6235 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][1] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n61 ) );
  INVX1 U6236 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n61 ), 
        .Y(n5607) );
  AND2X1 U6237 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][1] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n64 ) );
  INVX1 U6238 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n64 ), 
        .Y(n5608) );
  AND2X1 U6239 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][2] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n74 ) );
  INVX1 U6240 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n74 ), 
        .Y(n5609) );
  AND2X1 U6241 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][2] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n77 ) );
  INVX1 U6242 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n77 ), 
        .Y(n5610) );
  AND2X1 U6243 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][2] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n82 ) );
  INVX1 U6244 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n82 ), 
        .Y(n5611) );
  AND2X1 U6245 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][2] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n85 ) );
  INVX1 U6246 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n85 ), 
        .Y(n5612) );
  AND2X1 U6247 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][3] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n95 ) );
  INVX1 U6248 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n95 ), 
        .Y(n5613) );
  AND2X1 U6249 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][3] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n98 ) );
  INVX1 U6250 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n98 ), 
        .Y(n5614) );
  AND2X1 U6251 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][3] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n103 )
         );
  INVX1 U6252 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n103 ), 
        .Y(n5615) );
  AND2X1 U6253 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][3] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n106 )
         );
  INVX1 U6254 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n106 ), 
        .Y(n5616) );
  AND2X1 U6255 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][4] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n116 )
         );
  INVX1 U6256 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n116 ), 
        .Y(n5617) );
  AND2X1 U6257 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][4] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n119 )
         );
  INVX1 U6258 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n119 ), 
        .Y(n5618) );
  AND2X1 U6259 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][4] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n124 )
         );
  INVX1 U6260 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n124 ), 
        .Y(n5619) );
  AND2X1 U6261 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][4] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n127 )
         );
  INVX1 U6262 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n127 ), 
        .Y(n5620) );
  AND2X1 U6263 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][5] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n137 )
         );
  INVX1 U6264 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n137 ), 
        .Y(n5621) );
  AND2X1 U6265 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][5] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n140 )
         );
  INVX1 U6266 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n140 ), 
        .Y(n5622) );
  AND2X1 U6267 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][5] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n145 )
         );
  INVX1 U6268 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n145 ), 
        .Y(n5623) );
  AND2X1 U6269 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][5] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n148 )
         );
  INVX1 U6270 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n148 ), 
        .Y(n5624) );
  AND2X1 U6271 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][6] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n158 )
         );
  INVX1 U6272 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n158 ), 
        .Y(n5625) );
  AND2X1 U6273 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][6] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n161 )
         );
  INVX1 U6274 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n161 ), 
        .Y(n5626) );
  AND2X1 U6275 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][6] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n166 )
         );
  INVX1 U6276 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n166 ), 
        .Y(n5627) );
  AND2X1 U6277 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][6] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n169 )
         );
  INVX1 U6278 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n169 ), 
        .Y(n5628) );
  AND2X1 U6279 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][7] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n179 )
         );
  INVX1 U6280 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n179 ), 
        .Y(n5629) );
  AND2X1 U6281 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][7] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n182 )
         );
  INVX1 U6282 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n182 ), 
        .Y(n5630) );
  AND2X1 U6283 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][7] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n187 )
         );
  INVX1 U6284 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n187 ), 
        .Y(n5631) );
  AND2X1 U6285 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][7] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n190 )
         );
  INVX1 U6286 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n190 ), 
        .Y(n5632) );
  AND2X1 U6287 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][8] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n200 )
         );
  INVX1 U6288 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n200 ), 
        .Y(n5633) );
  AND2X1 U6289 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][8] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n203 )
         );
  INVX1 U6290 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n203 ), 
        .Y(n5634) );
  AND2X1 U6291 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][8] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n208 )
         );
  INVX1 U6292 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n208 ), 
        .Y(n5635) );
  AND2X1 U6293 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][8] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n211 )
         );
  INVX1 U6294 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n211 ), 
        .Y(n5636) );
  AND2X1 U6295 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][9] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n221 )
         );
  INVX1 U6296 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n221 ), 
        .Y(n5637) );
  AND2X1 U6297 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][9] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n224 )
         );
  INVX1 U6298 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n224 ), 
        .Y(n5638) );
  AND2X1 U6299 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][9] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n229 )
         );
  INVX1 U6300 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n229 ), 
        .Y(n5639) );
  AND2X1 U6301 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][9] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n232 )
         );
  INVX1 U6302 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n232 ), 
        .Y(n5640) );
  AND2X1 U6303 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][10] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n242 )
         );
  INVX1 U6304 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n242 ), 
        .Y(n5641) );
  AND2X1 U6305 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][10] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n245 )
         );
  INVX1 U6306 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n245 ), 
        .Y(n5642) );
  AND2X1 U6307 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][10] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n250 )
         );
  INVX1 U6308 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n250 ), 
        .Y(n5643) );
  AND2X1 U6309 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][10] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n253 )
         );
  INVX1 U6310 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n253 ), 
        .Y(n5644) );
  AND2X1 U6311 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][11] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n263 )
         );
  INVX1 U6312 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n263 ), 
        .Y(n5645) );
  AND2X1 U6313 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][11] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n266 )
         );
  INVX1 U6314 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n266 ), 
        .Y(n5646) );
  AND2X1 U6315 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][11] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n271 )
         );
  INVX1 U6316 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n271 ), 
        .Y(n5647) );
  AND2X1 U6317 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][11] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n274 )
         );
  INVX1 U6318 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n274 ), 
        .Y(n5648) );
  AND2X1 U6319 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][12] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n284 )
         );
  INVX1 U6320 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n284 ), 
        .Y(n5649) );
  AND2X1 U6321 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][12] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n287 )
         );
  INVX1 U6322 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n287 ), 
        .Y(n5650) );
  AND2X1 U6323 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][12] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n292 )
         );
  INVX1 U6324 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n292 ), 
        .Y(n5651) );
  AND2X1 U6325 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][12] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n295 )
         );
  INVX1 U6326 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n295 ), 
        .Y(n5652) );
  AND2X1 U6327 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][13] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n305 )
         );
  INVX1 U6328 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n305 ), 
        .Y(n5653) );
  AND2X1 U6329 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][13] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n308 )
         );
  INVX1 U6330 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n308 ), 
        .Y(n5654) );
  AND2X1 U6331 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][13] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n313 )
         );
  INVX1 U6332 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n313 ), 
        .Y(n5655) );
  AND2X1 U6333 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][13] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n316 )
         );
  INVX1 U6334 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n316 ), 
        .Y(n5656) );
  AND2X1 U6335 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][14] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n326 )
         );
  INVX1 U6336 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n326 ), 
        .Y(n5657) );
  AND2X1 U6337 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][14] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n329 )
         );
  INVX1 U6338 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n329 ), 
        .Y(n5658) );
  AND2X1 U6339 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][14] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n334 )
         );
  INVX1 U6340 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n334 ), 
        .Y(n5659) );
  AND2X1 U6341 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][14] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n337 )
         );
  INVX1 U6342 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n337 ), 
        .Y(n5660) );
  AND2X1 U6343 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][15] ), .B(n8878), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n347 )
         );
  INVX1 U6344 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n347 ), 
        .Y(n5661) );
  AND2X1 U6345 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][15] ), .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n350 )
         );
  INVX1 U6346 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n350 ), 
        .Y(n5662) );
  AND2X1 U6347 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][15] ), .B(n9821), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n358 )
         );
  INVX1 U6348 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n358 ), 
        .Y(n5663) );
  AND2X1 U6349 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][15] ), .B(n9817), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n368 )
         );
  INVX1 U6350 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n368 ), 
        .Y(n5664) );
  AND2X1 U6351 ( .A(a_length[31]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n153 ) );
  INVX1 U6352 ( .A(\Decision_AXILiteS_s_axi_U/n153 ), .Y(n5665) );
  AND2X1 U6353 ( .A(a_length[30]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n161 ) );
  INVX1 U6354 ( .A(\Decision_AXILiteS_s_axi_U/n161 ), .Y(n5666) );
  AND2X1 U6355 ( .A(a_length[29]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n164 ) );
  INVX1 U6356 ( .A(\Decision_AXILiteS_s_axi_U/n164 ), .Y(n5667) );
  AND2X1 U6357 ( .A(a_length[28]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n167 ) );
  INVX1 U6358 ( .A(\Decision_AXILiteS_s_axi_U/n167 ), .Y(n5668) );
  AND2X1 U6359 ( .A(a_length[27]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n170 ) );
  INVX1 U6360 ( .A(\Decision_AXILiteS_s_axi_U/n170 ), .Y(n5669) );
  AND2X1 U6361 ( .A(a_length[26]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n173 ) );
  INVX1 U6362 ( .A(\Decision_AXILiteS_s_axi_U/n173 ), .Y(n5670) );
  AND2X1 U6363 ( .A(a_length[25]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n176 ) );
  INVX1 U6364 ( .A(\Decision_AXILiteS_s_axi_U/n176 ), .Y(n5671) );
  AND2X1 U6365 ( .A(a_length[24]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n179 ) );
  INVX1 U6366 ( .A(\Decision_AXILiteS_s_axi_U/n179 ), .Y(n5672) );
  AND2X1 U6367 ( .A(a_length[23]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n182 ) );
  INVX1 U6368 ( .A(\Decision_AXILiteS_s_axi_U/n182 ), .Y(n5673) );
  AND2X1 U6369 ( .A(a_length[22]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n185 ) );
  INVX1 U6370 ( .A(\Decision_AXILiteS_s_axi_U/n185 ), .Y(n5674) );
  AND2X1 U6371 ( .A(a_length[21]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n188 ) );
  INVX1 U6372 ( .A(\Decision_AXILiteS_s_axi_U/n188 ), .Y(n5675) );
  AND2X1 U6373 ( .A(a_length[20]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n191 ) );
  INVX1 U6374 ( .A(\Decision_AXILiteS_s_axi_U/n191 ), .Y(n5676) );
  AND2X1 U6375 ( .A(a_length[19]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n194 ) );
  INVX1 U6376 ( .A(\Decision_AXILiteS_s_axi_U/n194 ), .Y(n5677) );
  AND2X1 U6377 ( .A(a_length[18]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n197 ) );
  INVX1 U6378 ( .A(\Decision_AXILiteS_s_axi_U/n197 ), .Y(n5678) );
  AND2X1 U6379 ( .A(a_length[17]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n200 ) );
  INVX1 U6380 ( .A(\Decision_AXILiteS_s_axi_U/n200 ), .Y(n5679) );
  AND2X1 U6381 ( .A(a_length[16]), .B(\Decision_AXILiteS_s_axi_U/n157 ), .Y(
        \Decision_AXILiteS_s_axi_U/n203 ) );
  INVX1 U6382 ( .A(\Decision_AXILiteS_s_axi_U/n203 ), .Y(n5680) );
  AND2X1 U6383 ( .A(s_axi_AXILiteS_RDATA[15]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n206 ) );
  INVX1 U6384 ( .A(\Decision_AXILiteS_s_axi_U/n206 ), .Y(n5681) );
  AND2X1 U6385 ( .A(s_axi_AXILiteS_RDATA[14]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n213 ) );
  INVX1 U6386 ( .A(\Decision_AXILiteS_s_axi_U/n213 ), .Y(n5682) );
  AND2X1 U6387 ( .A(s_axi_AXILiteS_RDATA[13]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n218 ) );
  INVX1 U6388 ( .A(\Decision_AXILiteS_s_axi_U/n218 ), .Y(n5683) );
  AND2X1 U6389 ( .A(s_axi_AXILiteS_RDATA[12]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n223 ) );
  INVX1 U6390 ( .A(\Decision_AXILiteS_s_axi_U/n223 ), .Y(n5684) );
  AND2X1 U6391 ( .A(s_axi_AXILiteS_RDATA[11]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n228 ) );
  INVX1 U6392 ( .A(\Decision_AXILiteS_s_axi_U/n228 ), .Y(n5685) );
  AND2X1 U6393 ( .A(s_axi_AXILiteS_RDATA[10]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n233 ) );
  INVX1 U6394 ( .A(\Decision_AXILiteS_s_axi_U/n233 ), .Y(n5686) );
  AND2X1 U6395 ( .A(s_axi_AXILiteS_RDATA[9]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n238 ) );
  INVX1 U6396 ( .A(\Decision_AXILiteS_s_axi_U/n238 ), .Y(n5687) );
  AND2X1 U6397 ( .A(s_axi_AXILiteS_RDATA[8]), .B(n8918), .Y(
        \Decision_AXILiteS_s_axi_U/n243 ) );
  INVX1 U6398 ( .A(\Decision_AXILiteS_s_axi_U/n243 ), .Y(n5688) );
  AND2X1 U6399 ( .A(vthresh[7]), .B(n9310), .Y(
        \Decision_AXILiteS_s_axi_U/n256 ) );
  INVX1 U6400 ( .A(\Decision_AXILiteS_s_axi_U/n256 ), .Y(n5689) );
  AND2X1 U6401 ( .A(vthresh[3]), .B(n9310), .Y(
        \Decision_AXILiteS_s_axi_U/n286 ) );
  INVX1 U6402 ( .A(\Decision_AXILiteS_s_axi_U/n286 ), .Y(n5690) );
  AND2X1 U6403 ( .A(vthresh[2]), .B(n9310), .Y(
        \Decision_AXILiteS_s_axi_U/n295 ) );
  INVX1 U6404 ( .A(\Decision_AXILiteS_s_axi_U/n295 ), .Y(n5691) );
  AND2X1 U6405 ( .A(athresh[1]), .B(n9309), .Y(
        \Decision_AXILiteS_s_axi_U/n305 ) );
  INVX1 U6406 ( .A(\Decision_AXILiteS_s_axi_U/n305 ), .Y(n5692) );
  AND2X1 U6407 ( .A(a_length[0]), .B(n9312), .Y(
        \Decision_AXILiteS_s_axi_U/n327 ) );
  INVX1 U6408 ( .A(\Decision_AXILiteS_s_axi_U/n327 ), .Y(n5693) );
  AND2X1 U6409 ( .A(n9900), .B(n349), .Y(n362) );
  INVX1 U6410 ( .A(n362), .Y(n5694) );
  AND2X1 U6411 ( .A(i_fu_607_p2[1]), .B(n349), .Y(n359) );
  INVX1 U6412 ( .A(n359), .Y(n5695) );
  BUFX2 U6413 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n12 ), 
        .Y(n5696) );
  BUFX2 U6414 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n7 ), 
        .Y(n5697) );
  BUFX2 U6415 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n12 ), 
        .Y(n5698) );
  BUFX2 U6416 ( .A(\Decision_AXILiteS_s_axi_U/n330 ), .Y(n5699) );
  BUFX2 U6417 ( .A(n11173), .Y(n5700) );
  BUFX2 U6418 ( .A(n11550), .Y(n5701) );
  BUFX2 U6419 ( .A(n11630), .Y(n5702) );
  BUFX2 U6420 ( .A(n11627), .Y(n5703) );
  BUFX2 U6421 ( .A(n11719), .Y(n5704) );
  BUFX2 U6422 ( .A(n11808), .Y(n5705) );
  BUFX2 U6423 ( .A(n11897), .Y(n5706) );
  BUFX2 U6424 ( .A(n12005), .Y(n5707) );
  BUFX2 U6425 ( .A(n12094), .Y(n5708) );
  BUFX2 U6426 ( .A(n12183), .Y(n5709) );
  BUFX2 U6427 ( .A(n12263), .Y(n5710) );
  BUFX2 U6428 ( .A(n12260), .Y(n5711) );
  INVX1 U6429 ( .A(\Decision_AXILiteS_s_axi_U/n301 ), .Y(n5713) );
  INVX1 U6430 ( .A(\Decision_AXILiteS_s_axi_U/n316 ), .Y(n5716) );
  BUFX2 U6431 ( .A(n1650), .Y(n5718) );
  INVX1 U6432 ( .A(\Decision_AXILiteS_s_axi_U/n252 ), .Y(n5719) );
  INVX1 U6433 ( .A(\Decision_AXILiteS_s_axi_U/n282 ), .Y(n5720) );
  INVX1 U6434 ( .A(\Decision_AXILiteS_s_axi_U/n291 ), .Y(n5721) );
  BUFX2 U6435 ( .A(n11497), .Y(n5722) );
  BUFX2 U6436 ( .A(n11534), .Y(n5723) );
  BUFX2 U6437 ( .A(n11541), .Y(n5724) );
  BUFX2 U6438 ( .A(n11666), .Y(n5725) );
  BUFX2 U6439 ( .A(n11703), .Y(n5726) );
  BUFX2 U6440 ( .A(n11710), .Y(n5727) );
  BUFX2 U6441 ( .A(n11755), .Y(n5728) );
  BUFX2 U6442 ( .A(n11792), .Y(n5729) );
  BUFX2 U6443 ( .A(n11799), .Y(n5730) );
  BUFX2 U6444 ( .A(n11989), .Y(n5731) );
  BUFX2 U6445 ( .A(n11996), .Y(n5732) );
  BUFX2 U6446 ( .A(n12085), .Y(n5733) );
  BUFX2 U6447 ( .A(n12130), .Y(n5734) );
  BUFX2 U6448 ( .A(n12167), .Y(n5735) );
  BUFX2 U6449 ( .A(n12174), .Y(n5736) );
  BUFX2 U6450 ( .A(n11065), .Y(n5737) );
  BUFX2 U6451 ( .A(n11083), .Y(n5738) );
  BUFX2 U6452 ( .A(n11125), .Y(n5739) );
  BUFX2 U6453 ( .A(n11485), .Y(n5740) );
  BUFX2 U6454 ( .A(n11502), .Y(n5741) );
  BUFX2 U6455 ( .A(n11565), .Y(n5742) );
  BUFX2 U6456 ( .A(n11654), .Y(n5743) );
  BUFX2 U6457 ( .A(n11671), .Y(n5744) );
  BUFX2 U6458 ( .A(n11743), .Y(n5745) );
  BUFX2 U6459 ( .A(n11760), .Y(n5746) );
  BUFX2 U6460 ( .A(n11849), .Y(n5747) );
  BUFX2 U6461 ( .A(n11940), .Y(n5748) );
  BUFX2 U6462 ( .A(n11957), .Y(n5749) );
  BUFX2 U6463 ( .A(n12046), .Y(n5750) );
  BUFX2 U6464 ( .A(n12118), .Y(n5751) );
  BUFX2 U6465 ( .A(n12135), .Y(n5752) );
  BUFX2 U6466 ( .A(n12198), .Y(n5753) );
  OR2X1 U6467 ( .A(n11059), .B(n7834), .Y(n11060) );
  INVX1 U6468 ( .A(n11060), .Y(n5754) );
  BUFX2 U6469 ( .A(n11064), .Y(n5755) );
  BUFX2 U6470 ( .A(n11082), .Y(n5756) );
  BUFX2 U6471 ( .A(n11061), .Y(n5757) );
  BUFX2 U6472 ( .A(n11080), .Y(n5758) );
  BUFX2 U6473 ( .A(n11127), .Y(n5759) );
  BUFX2 U6474 ( .A(n11504), .Y(n5760) );
  BUFX2 U6475 ( .A(n11610), .Y(n5761) );
  BUFX2 U6476 ( .A(n11624), .Y(n5762) );
  BUFX2 U6477 ( .A(n11673), .Y(n5763) );
  BUFX2 U6478 ( .A(n11762), .Y(n5764) );
  BUFX2 U6479 ( .A(n11851), .Y(n5765) );
  BUFX2 U6480 ( .A(n11959), .Y(n5766) );
  BUFX2 U6481 ( .A(n12048), .Y(n5767) );
  BUFX2 U6482 ( .A(n12137), .Y(n5768) );
  BUFX2 U6483 ( .A(n12243), .Y(n5769) );
  BUFX2 U6484 ( .A(n12257), .Y(n5770) );
  BUFX2 U6485 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n12 ), 
        .Y(n5771) );
  BUFX2 U6486 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n20 ), 
        .Y(n5772) );
  BUFX2 U6487 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n30 ), 
        .Y(n5773) );
  BUFX2 U6488 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n38 ), 
        .Y(n5774) );
  BUFX2 U6489 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n54 ), 
        .Y(n5775) );
  BUFX2 U6490 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n57 ), 
        .Y(n5776) );
  BUFX2 U6491 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n62 ), 
        .Y(n5777) );
  BUFX2 U6492 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n65 ), 
        .Y(n5778) );
  BUFX2 U6493 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n75 ), 
        .Y(n5779) );
  BUFX2 U6494 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n78 ), 
        .Y(n5780) );
  BUFX2 U6495 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n83 ), 
        .Y(n5781) );
  BUFX2 U6496 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n86 ), 
        .Y(n5782) );
  BUFX2 U6497 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n96 ), 
        .Y(n5783) );
  BUFX2 U6498 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n99 ), 
        .Y(n5784) );
  BUFX2 U6499 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n104 ), 
        .Y(n5785) );
  BUFX2 U6500 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n107 ), 
        .Y(n5786) );
  BUFX2 U6501 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n117 ), 
        .Y(n5787) );
  BUFX2 U6502 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n120 ), 
        .Y(n5788) );
  BUFX2 U6503 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n125 ), 
        .Y(n5789) );
  BUFX2 U6504 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n128 ), 
        .Y(n5790) );
  BUFX2 U6505 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n138 ), 
        .Y(n5791) );
  BUFX2 U6506 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n141 ), 
        .Y(n5792) );
  BUFX2 U6507 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n146 ), 
        .Y(n5793) );
  BUFX2 U6508 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n149 ), 
        .Y(n5794) );
  BUFX2 U6509 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n159 ), 
        .Y(n5795) );
  BUFX2 U6510 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n162 ), 
        .Y(n5796) );
  BUFX2 U6511 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n167 ), 
        .Y(n5797) );
  BUFX2 U6512 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n170 ), 
        .Y(n5798) );
  BUFX2 U6513 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n180 ), 
        .Y(n5799) );
  BUFX2 U6514 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n183 ), 
        .Y(n5800) );
  BUFX2 U6515 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n188 ), 
        .Y(n5801) );
  BUFX2 U6516 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n191 ), 
        .Y(n5802) );
  BUFX2 U6517 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n201 ), 
        .Y(n5803) );
  BUFX2 U6518 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n204 ), 
        .Y(n5804) );
  BUFX2 U6519 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n209 ), 
        .Y(n5805) );
  BUFX2 U6520 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n212 ), 
        .Y(n5806) );
  BUFX2 U6521 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n222 ), 
        .Y(n5807) );
  BUFX2 U6522 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n225 ), 
        .Y(n5808) );
  BUFX2 U6523 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n230 ), 
        .Y(n5809) );
  BUFX2 U6524 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n233 ), 
        .Y(n5810) );
  BUFX2 U6525 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n243 ), 
        .Y(n5811) );
  BUFX2 U6526 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n246 ), 
        .Y(n5812) );
  BUFX2 U6527 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n251 ), 
        .Y(n5813) );
  BUFX2 U6528 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n254 ), 
        .Y(n5814) );
  BUFX2 U6529 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n264 ), 
        .Y(n5815) );
  BUFX2 U6530 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n267 ), 
        .Y(n5816) );
  BUFX2 U6531 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n272 ), 
        .Y(n5817) );
  BUFX2 U6532 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n275 ), 
        .Y(n5818) );
  BUFX2 U6533 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n285 ), 
        .Y(n5819) );
  BUFX2 U6534 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n288 ), 
        .Y(n5820) );
  BUFX2 U6535 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n293 ), 
        .Y(n5821) );
  BUFX2 U6536 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n296 ), 
        .Y(n5822) );
  BUFX2 U6537 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n306 ), 
        .Y(n5823) );
  BUFX2 U6538 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n309 ), 
        .Y(n5824) );
  BUFX2 U6539 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n314 ), 
        .Y(n5825) );
  BUFX2 U6540 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n317 ), 
        .Y(n5826) );
  BUFX2 U6541 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n327 ), 
        .Y(n5827) );
  BUFX2 U6542 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n330 ), 
        .Y(n5828) );
  BUFX2 U6543 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n335 ), 
        .Y(n5829) );
  BUFX2 U6544 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n338 ), 
        .Y(n5830) );
  BUFX2 U6545 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n348 ), 
        .Y(n5831) );
  BUFX2 U6546 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n351 ), 
        .Y(n5832) );
  BUFX2 U6547 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n359 ), 
        .Y(n5833) );
  BUFX2 U6548 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n369 ), 
        .Y(n5834) );
  BUFX2 U6549 ( .A(\Decision_AXILiteS_s_axi_U/n154 ), .Y(n5835) );
  BUFX2 U6550 ( .A(\Decision_AXILiteS_s_axi_U/n162 ), .Y(n5836) );
  BUFX2 U6551 ( .A(\Decision_AXILiteS_s_axi_U/n165 ), .Y(n5837) );
  BUFX2 U6552 ( .A(\Decision_AXILiteS_s_axi_U/n168 ), .Y(n5838) );
  BUFX2 U6553 ( .A(\Decision_AXILiteS_s_axi_U/n171 ), .Y(n5839) );
  BUFX2 U6554 ( .A(\Decision_AXILiteS_s_axi_U/n174 ), .Y(n5840) );
  BUFX2 U6555 ( .A(\Decision_AXILiteS_s_axi_U/n177 ), .Y(n5841) );
  BUFX2 U6556 ( .A(\Decision_AXILiteS_s_axi_U/n180 ), .Y(n5842) );
  BUFX2 U6557 ( .A(\Decision_AXILiteS_s_axi_U/n183 ), .Y(n5843) );
  BUFX2 U6558 ( .A(\Decision_AXILiteS_s_axi_U/n186 ), .Y(n5844) );
  BUFX2 U6559 ( .A(\Decision_AXILiteS_s_axi_U/n189 ), .Y(n5845) );
  BUFX2 U6560 ( .A(\Decision_AXILiteS_s_axi_U/n192 ), .Y(n5846) );
  BUFX2 U6561 ( .A(\Decision_AXILiteS_s_axi_U/n195 ), .Y(n5847) );
  BUFX2 U6562 ( .A(\Decision_AXILiteS_s_axi_U/n198 ), .Y(n5848) );
  BUFX2 U6563 ( .A(\Decision_AXILiteS_s_axi_U/n201 ), .Y(n5849) );
  BUFX2 U6564 ( .A(\Decision_AXILiteS_s_axi_U/n204 ), .Y(n5850) );
  BUFX2 U6565 ( .A(\Decision_AXILiteS_s_axi_U/n257 ), .Y(n5851) );
  BUFX2 U6566 ( .A(\Decision_AXILiteS_s_axi_U/n287 ), .Y(n5852) );
  BUFX2 U6567 ( .A(\Decision_AXILiteS_s_axi_U/n296 ), .Y(n5853) );
  INVX1 U6568 ( .A(n5855), .Y(n5854) );
  BUFX2 U6569 ( .A(\Decision_AXILiteS_s_axi_U/n303 ), .Y(n5855) );
  BUFX2 U6570 ( .A(\Decision_AXILiteS_s_axi_U/n306 ), .Y(n5856) );
  INVX1 U6571 ( .A(n5858), .Y(n5857) );
  BUFX2 U6572 ( .A(\Decision_AXILiteS_s_axi_U/n318 ), .Y(n5858) );
  BUFX2 U6573 ( .A(n363), .Y(n5859) );
  BUFX2 U6574 ( .A(n360), .Y(n5860) );
  BUFX2 U6575 ( .A(n11107), .Y(n5861) );
  BUFX2 U6576 ( .A(n11484), .Y(n5862) );
  BUFX2 U6577 ( .A(n11572), .Y(n5863) );
  BUFX2 U6578 ( .A(n11604), .Y(n5864) );
  BUFX2 U6579 ( .A(n11608), .Y(n5865) );
  BUFX2 U6580 ( .A(n11653), .Y(n5866) );
  BUFX2 U6581 ( .A(n11742), .Y(n5867) );
  BUFX2 U6582 ( .A(n11831), .Y(n5868) );
  BUFX2 U6583 ( .A(n11939), .Y(n5869) );
  BUFX2 U6584 ( .A(n12028), .Y(n5870) );
  BUFX2 U6585 ( .A(n12117), .Y(n5871) );
  BUFX2 U6586 ( .A(n12205), .Y(n5872) );
  BUFX2 U6587 ( .A(n12237), .Y(n5873) );
  BUFX2 U6588 ( .A(n12241), .Y(n5874) );
  BUFX2 U6589 ( .A(\Decision_AXILiteS_s_axi_U/n328 ), .Y(n5875) );
  AND2X1 U6590 ( .A(n11917), .B(n7587), .Y(N500) );
  INVX1 U6591 ( .A(N500), .Y(n5876) );
  AND2X1 U6592 ( .A(recentdatapoints_data_q0[0]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n3 ) );
  INVX1 U6593 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n3 ), 
        .Y(n5877) );
  AND2X1 U6594 ( .A(recentdatapoints_data_q0[1]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n47 ) );
  INVX1 U6595 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n47 ), 
        .Y(n5878) );
  AND2X1 U6596 ( .A(recentdatapoints_data_q0[2]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n68 ) );
  INVX1 U6597 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n68 ), 
        .Y(n5879) );
  AND2X1 U6598 ( .A(recentdatapoints_data_q0[3]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n89 ) );
  INVX1 U6599 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n89 ), 
        .Y(n5880) );
  AND2X1 U6600 ( .A(recentdatapoints_data_q0[4]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n110 )
         );
  INVX1 U6601 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n110 ), 
        .Y(n5881) );
  AND2X1 U6602 ( .A(recentdatapoints_data_q0[5]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n131 )
         );
  INVX1 U6603 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n131 ), 
        .Y(n5882) );
  AND2X1 U6604 ( .A(recentdatapoints_data_q0[6]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n152 )
         );
  INVX1 U6605 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n152 ), 
        .Y(n5883) );
  AND2X1 U6606 ( .A(recentdatapoints_data_q0[7]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n173 )
         );
  INVX1 U6607 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n173 ), 
        .Y(n5884) );
  AND2X1 U6608 ( .A(recentdatapoints_data_q0[8]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n194 )
         );
  INVX1 U6609 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n194 ), 
        .Y(n5885) );
  AND2X1 U6610 ( .A(recentdatapoints_data_q0[9]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n215 )
         );
  INVX1 U6611 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n215 ), 
        .Y(n5886) );
  AND2X1 U6612 ( .A(recentdatapoints_data_q0[10]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n236 )
         );
  INVX1 U6613 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n236 ), 
        .Y(n5887) );
  AND2X1 U6614 ( .A(recentdatapoints_data_q0[11]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n257 )
         );
  INVX1 U6615 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n257 ), 
        .Y(n5888) );
  AND2X1 U6616 ( .A(recentdatapoints_data_q0[12]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n278 )
         );
  INVX1 U6617 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n278 ), 
        .Y(n5889) );
  AND2X1 U6618 ( .A(recentdatapoints_data_q0[13]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n299 )
         );
  INVX1 U6619 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n299 ), 
        .Y(n5890) );
  AND2X1 U6620 ( .A(recentdatapoints_data_q0[14]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n320 )
         );
  INVX1 U6621 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n320 ), 
        .Y(n5891) );
  AND2X1 U6622 ( .A(recentdatapoints_data_q0[15]), .B(N472), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n341 )
         );
  INVX1 U6623 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n341 ), 
        .Y(n5892) );
  AND2X1 U6624 ( .A(\Decision_AXILiteS_s_axi_U/int_isr[1] ), .B(
        \Decision_AXILiteS_s_axi_U/n598 ), .Y(\Decision_AXILiteS_s_axi_U/n597 ) );
  INVX1 U6625 ( .A(\Decision_AXILiteS_s_axi_U/n597 ), .Y(n5893) );
  OR2X1 U6626 ( .A(n8859), .B(n8858), .Y(\Decision_AXILiteS_s_axi_U/n632 ) );
  INVX1 U6627 ( .A(\Decision_AXILiteS_s_axi_U/n632 ), .Y(n5894) );
  BUFX2 U6628 ( .A(n1675), .Y(n5895) );
  BUFX2 U6629 ( .A(n288), .Y(n5896) );
  BUFX2 U6630 ( .A(n264), .Y(n5897) );
  AND2X1 U6631 ( .A(\Decision_AXILiteS_s_axi_U/n310 ), .B(n8858), .Y(
        \Decision_AXILiteS_s_axi_U/n308 ) );
  INVX1 U6632 ( .A(\Decision_AXILiteS_s_axi_U/n308 ), .Y(n5898) );
  BUFX2 U6633 ( .A(n1676), .Y(n5899) );
  BUFX2 U6634 ( .A(n289), .Y(n5900) );
  AND2X1 U6635 ( .A(n276), .B(n277), .Y(n265) );
  INVX1 U6636 ( .A(n265), .Y(n5901) );
  BUFX2 U6637 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n21 ), 
        .Y(n5902) );
  BUFX2 U6638 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n20 ), 
        .Y(n5903) );
  BUFX2 U6639 ( .A(\Decision_AXILiteS_s_axi_U/n309 ), .Y(n5904) );
  AND2X1 U6640 ( .A(n9927), .B(n9926), .Y(n1677) );
  INVX1 U6641 ( .A(n1677), .Y(n5905) );
  AND2X1 U6642 ( .A(n10689), .B(n10691), .Y(n290) );
  INVX1 U6643 ( .A(n290), .Y(n5906) );
  AND2X1 U6644 ( .A(n267), .B(n268), .Y(n266) );
  INVX1 U6645 ( .A(n266), .Y(n5907) );
  AND2X1 U6646 ( .A(n11199), .B(n7441), .Y(n11200) );
  INVX1 U6647 ( .A(n11200), .Y(n5908) );
  AND2X1 U6648 ( .A(n11200), .B(n7644), .Y(n11201) );
  INVX1 U6649 ( .A(n11201), .Y(n5909) );
  AND2X1 U6650 ( .A(n11204), .B(n7860), .Y(n11175) );
  INVX1 U6651 ( .A(n11175), .Y(n5910) );
  AND2X1 U6652 ( .A(n11176), .B(n7439), .Y(n11177) );
  INVX1 U6653 ( .A(n11177), .Y(n5911) );
  AND2X1 U6654 ( .A(n11177), .B(n7642), .Y(n11178) );
  INVX1 U6655 ( .A(n11178), .Y(n5912) );
  AND2X1 U6656 ( .A(n11180), .B(n6254), .Y(n11181) );
  INVX1 U6657 ( .A(n11181), .Y(n5913) );
  AND2X1 U6658 ( .A(n11181), .B(n6351), .Y(n11182) );
  INVX1 U6659 ( .A(n11182), .Y(n5914) );
  AND2X1 U6660 ( .A(n11182), .B(n7443), .Y(n11183) );
  INVX1 U6661 ( .A(n11183), .Y(n5915) );
  AND2X1 U6662 ( .A(n11183), .B(n7864), .Y(n11185) );
  INVX1 U6663 ( .A(n11185), .Y(n5916) );
  AND2X1 U6664 ( .A(n11185), .B(n6460), .Y(n11186) );
  INVX1 U6665 ( .A(n11186), .Y(n5917) );
  AND2X1 U6666 ( .A(n11186), .B(n7265), .Y(n11187) );
  INVX1 U6667 ( .A(n11187), .Y(n5918) );
  AND2X1 U6668 ( .A(n11187), .B(n7100), .Y(n11188) );
  INVX1 U6669 ( .A(n11188), .Y(n5919) );
  AND2X1 U6670 ( .A(n11189), .B(n6573), .Y(n11190) );
  INVX1 U6671 ( .A(n11190), .Y(n5920) );
  AND2X1 U6672 ( .A(n11190), .B(n6948), .Y(n11191) );
  INVX1 U6673 ( .A(n11191), .Y(n5921) );
  AND2X1 U6674 ( .A(n11191), .B(n6813), .Y(n11192) );
  INVX1 U6675 ( .A(n11192), .Y(n5922) );
  AND2X1 U6676 ( .A(n11192), .B(n7646), .Y(n11193) );
  INVX1 U6677 ( .A(n11193), .Y(n5923) );
  AND2X1 U6678 ( .A(n11193), .B(n6688), .Y(n11194) );
  INVX1 U6679 ( .A(n11194), .Y(n5924) );
  AND2X1 U6680 ( .A(n11229), .B(n7440), .Y(n11230) );
  INVX1 U6681 ( .A(n11230), .Y(n5925) );
  AND2X1 U6682 ( .A(n11230), .B(n7643), .Y(n11231) );
  INVX1 U6683 ( .A(n11231), .Y(n5926) );
  AND2X1 U6684 ( .A(n11234), .B(n7859), .Y(n11205) );
  INVX1 U6685 ( .A(n11205), .Y(n5927) );
  AND2X1 U6686 ( .A(n11206), .B(n7438), .Y(n11207) );
  INVX1 U6687 ( .A(n11207), .Y(n5928) );
  AND2X1 U6688 ( .A(n11207), .B(n7641), .Y(n11208) );
  INVX1 U6689 ( .A(n11208), .Y(n5929) );
  AND2X1 U6690 ( .A(n11210), .B(n6253), .Y(n11211) );
  INVX1 U6691 ( .A(n11211), .Y(n5930) );
  AND2X1 U6692 ( .A(n11211), .B(n6350), .Y(n11212) );
  INVX1 U6693 ( .A(n11212), .Y(n5931) );
  AND2X1 U6694 ( .A(n11212), .B(n7442), .Y(n11213) );
  INVX1 U6695 ( .A(n11213), .Y(n5932) );
  AND2X1 U6696 ( .A(n11213), .B(n7863), .Y(n11215) );
  INVX1 U6697 ( .A(n11215), .Y(n5933) );
  AND2X1 U6698 ( .A(n11215), .B(n6459), .Y(n11216) );
  INVX1 U6699 ( .A(n11216), .Y(n5934) );
  AND2X1 U6700 ( .A(n11216), .B(n7264), .Y(n11217) );
  INVX1 U6701 ( .A(n11217), .Y(n5935) );
  AND2X1 U6702 ( .A(n11217), .B(n7099), .Y(n11218) );
  INVX1 U6703 ( .A(n11218), .Y(n5936) );
  AND2X1 U6704 ( .A(n11219), .B(n6572), .Y(n11220) );
  INVX1 U6705 ( .A(n11220), .Y(n5937) );
  AND2X1 U6706 ( .A(n11220), .B(n6947), .Y(n11221) );
  INVX1 U6707 ( .A(n11221), .Y(n5938) );
  AND2X1 U6708 ( .A(n11221), .B(n6812), .Y(n11222) );
  INVX1 U6709 ( .A(n11222), .Y(n5939) );
  AND2X1 U6710 ( .A(n11222), .B(n7645), .Y(n11223) );
  INVX1 U6711 ( .A(n11223), .Y(n5940) );
  AND2X1 U6712 ( .A(n11223), .B(n6687), .Y(n11224) );
  INVX1 U6713 ( .A(n11224), .Y(n5941) );
  INVX1 U6714 ( .A(n11562), .Y(n5943) );
  INVX1 U6715 ( .A(n12195), .Y(n5946) );
  INVX1 U6716 ( .A(n5949), .Y(n5948) );
  BUFX2 U6717 ( .A(n585), .Y(n5949) );
  AND2X1 U6718 ( .A(\tmp_22_reg_1772[0] ), .B(n10673), .Y(n685) );
  INVX1 U6719 ( .A(n685), .Y(n5950) );
  INVX1 U6720 ( .A(n5952), .Y(n5951) );
  BUFX2 U6721 ( .A(n11651), .Y(n5952) );
  INVX1 U6722 ( .A(n5954), .Y(n5953) );
  BUFX2 U6723 ( .A(n12115), .Y(n5954) );
  AND2X1 U6724 ( .A(s_axi_AXILiteS_WSTRB[0]), .B(ap_rst_n), .Y(
        \Decision_AXILiteS_s_axi_U/n617 ) );
  INVX1 U6725 ( .A(\Decision_AXILiteS_s_axi_U/n617 ), .Y(n5955) );
  INVX1 U6726 ( .A(n8372), .Y(n5957) );
  INVX1 U6727 ( .A(n8371), .Y(n5960) );
  BUFX2 U6728 ( .A(\Decision_AXILiteS_s_axi_U/n522 ), .Y(n5962) );
  INVX1 U6729 ( .A(n5964), .Y(n5963) );
  BUFX2 U6730 ( .A(\Decision_AXILiteS_s_axi_U/n622 ), .Y(n5964) );
  INVX1 U6731 ( .A(n5966), .Y(n5965) );
  BUFX2 U6732 ( .A(n2237), .Y(n5966) );
  AND2X1 U6733 ( .A(ACaptureThresh_loc_reg_288[19]), .B(n7864), .Y(n11698) );
  INVX1 U6734 ( .A(n11698), .Y(n5967) );
  AND2X1 U6735 ( .A(ACaptureThresh_loc_reg_288[27]), .B(n7646), .Y(n11681) );
  INVX1 U6736 ( .A(n11681), .Y(n5968) );
  AND2X1 U6737 ( .A(VCaptureThresh_loc_reg_298[19]), .B(n7863), .Y(n12162) );
  INVX1 U6738 ( .A(n12162), .Y(n5969) );
  AND2X1 U6739 ( .A(VCaptureThresh_loc_reg_298[27]), .B(n7645), .Y(n12145) );
  INVX1 U6740 ( .A(n12145), .Y(n5970) );
  INVX1 U6741 ( .A(n347), .Y(n5972) );
  INVX1 U6742 ( .A(n345), .Y(n5973) );
  BUFX2 U6743 ( .A(n11268), .Y(n5975) );
  BUFX2 U6744 ( .A(n11272), .Y(n5976) );
  BUFX2 U6745 ( .A(n11276), .Y(n5977) );
  BUFX2 U6746 ( .A(n11280), .Y(n5978) );
  BUFX2 U6747 ( .A(n11284), .Y(n5979) );
  BUFX2 U6748 ( .A(n11288), .Y(n5980) );
  BUFX2 U6749 ( .A(n11292), .Y(n5981) );
  BUFX2 U6750 ( .A(n11296), .Y(n5982) );
  BUFX2 U6751 ( .A(n11300), .Y(n5983) );
  BUFX2 U6752 ( .A(n11320), .Y(n5984) );
  BUFX2 U6753 ( .A(n11324), .Y(n5985) );
  BUFX2 U6754 ( .A(n11328), .Y(n5986) );
  BUFX2 U6755 ( .A(n11332), .Y(n5987) );
  BUFX2 U6756 ( .A(n11336), .Y(n5988) );
  BUFX2 U6757 ( .A(n11340), .Y(n5989) );
  BUFX2 U6758 ( .A(n11344), .Y(n5990) );
  BUFX2 U6759 ( .A(n11348), .Y(n5991) );
  BUFX2 U6760 ( .A(n11372), .Y(n5992) );
  BUFX2 U6761 ( .A(n11376), .Y(n5993) );
  BUFX2 U6762 ( .A(n11380), .Y(n5994) );
  BUFX2 U6763 ( .A(n11384), .Y(n5995) );
  BUFX2 U6764 ( .A(n11388), .Y(n5996) );
  BUFX2 U6765 ( .A(n11392), .Y(n5997) );
  BUFX2 U6766 ( .A(n11396), .Y(n5998) );
  BUFX2 U6767 ( .A(n11400), .Y(n5999) );
  BUFX2 U6768 ( .A(n11404), .Y(n6000) );
  BUFX2 U6769 ( .A(n11424), .Y(n6001) );
  BUFX2 U6770 ( .A(n11428), .Y(n6002) );
  BUFX2 U6771 ( .A(n11432), .Y(n6003) );
  BUFX2 U6772 ( .A(n11436), .Y(n6004) );
  BUFX2 U6773 ( .A(n11440), .Y(n6005) );
  BUFX2 U6774 ( .A(n11444), .Y(n6006) );
  BUFX2 U6775 ( .A(n11448), .Y(n6007) );
  BUFX2 U6776 ( .A(n11452), .Y(n6008) );
  INVX1 U6777 ( .A(\Decision_AXILiteS_s_axi_U/n612 ), .Y(n6009) );
  BUFX2 U6778 ( .A(n11697), .Y(n6010) );
  BUFX2 U6779 ( .A(n12161), .Y(n6011) );
  INVX1 U6780 ( .A(n357), .Y(n6013) );
  INVX1 U6781 ( .A(n355), .Y(n6014) );
  INVX1 U6782 ( .A(recentABools_data_address0[4]), .Y(n6016) );
  INVX1 U6783 ( .A(recentVBools_data_address0[4]), .Y(n6017) );
  BUFX2 U6784 ( .A(n6019), .Y(n6018) );
  INVX1 U6785 ( .A(n354), .Y(n6020) );
  INVX1 U6786 ( .A(n352), .Y(n6021) );
  AND2X1 U6787 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n73 ), .B(recentABools_data_address0[0]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n48 ) );
  INVX1 U6788 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n48 ), 
        .Y(n6023) );
  INVX1 U6789 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n19 ), 
        .Y(n6025) );
  AND2X1 U6790 ( .A(n9019), .B(n8049), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n19 ) );
  INVX1 U6791 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n18 ), 
        .Y(n6028) );
  AND2X1 U6792 ( .A(ap_CS_fsm[4]), .B(n7825), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n18 ) );
  BUFX2 U6793 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n44 ), 
        .Y(n6030) );
  BUFX2 U6794 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n46 ), 
        .Y(n6031) );
  AND2X1 U6795 ( .A(n10059), .B(\tmp_12_reg_1694[0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n53 ) );
  INVX1 U6796 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n53 ), 
        .Y(n6032) );
  AND2X1 U6797 ( .A(n10058), .B(\tmp_12_reg_1694[0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n64 ) );
  INVX1 U6798 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n64 ), 
        .Y(n6033) );
  AND2X1 U6799 ( .A(n9931), .B(\tmp_s_reg_1578[0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n51 ) );
  INVX1 U6800 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n51 ), 
        .Y(n6034) );
  AND2X1 U6801 ( .A(n9930), .B(\tmp_s_reg_1578[0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n62 ) );
  INVX1 U6802 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n62 ), 
        .Y(n6035) );
  AND2X1 U6803 ( .A(a_length[4]), .B(n8952), .Y(n3118) );
  INVX1 U6804 ( .A(n3118), .Y(n6036) );
  AND2X1 U6805 ( .A(a_length[17]), .B(n8953), .Y(n3092) );
  INVX1 U6806 ( .A(n3092), .Y(n6037) );
  AND2X1 U6807 ( .A(v_length[1]), .B(n8954), .Y(n2996) );
  INVX1 U6808 ( .A(n2996), .Y(n6038) );
  AND2X1 U6809 ( .A(recentdatapoints_head_i[9]), .B(n8980), .Y(n1974) );
  INVX1 U6810 ( .A(n1974), .Y(n6039) );
  AND2X1 U6811 ( .A(recentdatapoints_head_i[19]), .B(n8979), .Y(n1964) );
  INVX1 U6812 ( .A(n1964), .Y(n6040) );
  AND2X1 U6813 ( .A(recentVBools_head_i[5]), .B(n9011), .Y(n1789) );
  INVX1 U6814 ( .A(n1789), .Y(n6041) );
  AND2X1 U6815 ( .A(recentVBools_head_i[12]), .B(n9010), .Y(n1768) );
  INVX1 U6816 ( .A(n1768), .Y(n6042) );
  AND2X1 U6817 ( .A(recentVBools_head_i[19]), .B(n9009), .Y(n1747) );
  INVX1 U6818 ( .A(n1747), .Y(n6043) );
  AND2X1 U6819 ( .A(CircularBuffer_head_i_read_ass_reg_1624[29]), .B(n9008), 
        .Y(n1718) );
  INVX1 U6820 ( .A(n1718), .Y(n6044) );
  AND2X1 U6821 ( .A(n2772), .B(n8992), .Y(n1631) );
  INVX1 U6822 ( .A(n1631), .Y(n6045) );
  AND2X1 U6823 ( .A(n2764), .B(n8993), .Y(n1625) );
  INVX1 U6824 ( .A(n1625), .Y(n6046) );
  BUFX2 U6825 ( .A(n2859), .Y(n6047) );
  BUFX2 U6826 ( .A(n2835), .Y(n6048) );
  AND2X1 U6827 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[2]), .Y(n2688) );
  INVX1 U6828 ( .A(n2688), .Y(n6049) );
  AND2X1 U6829 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[28]), .B(n9033), 
        .Y(n1396) );
  INVX1 U6830 ( .A(n1396), .Y(n6050) );
  AND2X1 U6831 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[6]), .B(n9036), 
        .Y(n1352) );
  INVX1 U6832 ( .A(n1352), .Y(n6051) );
  AND2X1 U6833 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[0]), .B(n9037), 
        .Y(n1334) );
  INVX1 U6834 ( .A(n1334), .Y(n6052) );
  AND2X1 U6835 ( .A(recentABools_head_i[6]), .B(n9038), .Y(n1329) );
  INVX1 U6836 ( .A(n1329), .Y(n6053) );
  AND2X1 U6837 ( .A(recentABools_head_i[9]), .B(n9039), .Y(n1322) );
  INVX1 U6838 ( .A(n1322), .Y(n6054) );
  AND2X1 U6839 ( .A(VbeatFallDelay_new_1_reg_342[0]), .B(n9013), .Y(n2157) );
  INVX1 U6840 ( .A(n2157), .Y(n6055) );
  AND2X1 U6841 ( .A(tmp_5_fu_726_p2[21]), .B(n8994), .Y(n1124) );
  INVX1 U6842 ( .A(n1124), .Y(n6056) );
  AND2X1 U6843 ( .A(tmp_4_fu_716_p2[8]), .B(n8995), .Y(n1053) );
  INVX1 U6844 ( .A(n1053), .Y(n6057) );
  AND2X1 U6845 ( .A(tmp_4_fu_716_p2[27]), .B(n8996), .Y(n989) );
  INVX1 U6846 ( .A(n989), .Y(n6058) );
  AND2X1 U6847 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[7]), .Y(n2434) );
  INVX1 U6848 ( .A(n2434), .Y(n6059) );
  AND2X1 U6849 ( .A(AbeatDelay[7]), .B(n10670), .Y(n767) );
  INVX1 U6850 ( .A(n767), .Y(n6060) );
  AND2X1 U6851 ( .A(tmp_3_fu_706_p2[14]), .B(n8997), .Y(n746) );
  INVX1 U6852 ( .A(n746), .Y(n6061) );
  AND2X1 U6853 ( .A(AbeatDelay[18]), .B(n8896), .Y(n730) );
  INVX1 U6854 ( .A(n730), .Y(n6062) );
  AND2X1 U6855 ( .A(AstimDelay[7]), .B(n8896), .Y(n662) );
  INVX1 U6856 ( .A(n662), .Y(n6063) );
  AND2X1 U6857 ( .A(tmp_6_fu_497_p3[11]), .B(n8966), .Y(n651) );
  INVX1 U6858 ( .A(n651), .Y(n6064) );
  AND2X1 U6859 ( .A(AstimDelay[24]), .B(n10670), .Y(n611) );
  INVX1 U6860 ( .A(n611), .Y(n6065) );
  AND2X1 U6861 ( .A(VstimDelay[10]), .B(n10670), .Y(n553) );
  INVX1 U6862 ( .A(n553), .Y(n6066) );
  AND2X1 U6863 ( .A(tmp_7_fu_511_p3[13]), .B(n8964), .Y(n545) );
  INVX1 U6864 ( .A(n545), .Y(n6067) );
  AND2X1 U6865 ( .A(\Decision_AXILiteS_s_axi_U/n564 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n416 ) );
  INVX1 U6866 ( .A(\Decision_AXILiteS_s_axi_U/n416 ), .Y(n6068) );
  AND2X1 U6867 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[2]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n383 )
         );
  INVX1 U6868 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n383 ), 
        .Y(n6069) );
  AND2X1 U6869 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[8]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n395 )
         );
  INVX1 U6870 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n395 ), 
        .Y(n6070) );
  AND2X1 U6871 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[7]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n428 )
         );
  INVX1 U6872 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n428 ), 
        .Y(n6071) );
  AND2X1 U6873 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[6]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n460 )
         );
  INVX1 U6874 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n460 ), 
        .Y(n6072) );
  AND2X1 U6875 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[1]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n484 )
         );
  INVX1 U6876 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n484 ), 
        .Y(n6073) );
  AND2X1 U6877 ( .A(n9467), .B(data_read_reg_1495[0]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n516 )
         );
  INVX1 U6878 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n516 ), 
        .Y(n6074) );
  AND2X1 U6879 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][10] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n571 )
         );
  INVX1 U6880 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n571 ), 
        .Y(n6075) );
  AND2X1 U6881 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][9] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n662 )
         );
  INVX1 U6882 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n662 ), 
        .Y(n6076) );
  AND2X1 U6883 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][8] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n680 )
         );
  INVX1 U6884 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n680 ), 
        .Y(n6077) );
  AND2X1 U6885 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][7] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n697 )
         );
  INVX1 U6886 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n697 ), 
        .Y(n6078) );
  AND2X1 U6887 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][6] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n713 )
         );
  INVX1 U6888 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n713 ), 
        .Y(n6079) );
  AND2X1 U6889 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][5] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n729 )
         );
  INVX1 U6890 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n729 ), 
        .Y(n6080) );
  AND2X1 U6891 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][4] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n745 )
         );
  INVX1 U6892 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n745 ), 
        .Y(n6081) );
  AND2X1 U6893 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][3] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n761 )
         );
  INVX1 U6894 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n761 ), 
        .Y(n6082) );
  AND2X1 U6895 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][2] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n811 )
         );
  INVX1 U6896 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n811 ), 
        .Y(n6083) );
  AND2X1 U6897 ( .A(sum_reg_308[7]), .B(n8929), .Y(n2670) );
  INVX1 U6898 ( .A(n2670), .Y(n6084) );
  AND2X1 U6899 ( .A(sum_1_reg_376[8]), .B(n8930), .Y(n2440) );
  INVX1 U6900 ( .A(n2440), .Y(n6085) );
  INVX1 U6901 ( .A(n4631), .Y(n6086) );
  AND2X1 U6902 ( .A(ACaptureThresh_loc_reg_288[3]), .B(n8968), .Y(n3056) );
  INVX1 U6903 ( .A(n3056), .Y(n6087) );
  BUFX2 U6904 ( .A(n3055), .Y(n6088) );
  BUFX2 U6905 ( .A(n3186), .Y(n6089) );
  BUFX2 U6906 ( .A(n3185), .Y(n6090) );
  BUFX2 U6907 ( .A(n3238), .Y(n6091) );
  BUFX2 U6908 ( .A(n3237), .Y(n6092) );
  AND2X1 U6909 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[1]), 
        .Y(n458) );
  INVX1 U6910 ( .A(n458), .Y(n6093) );
  BUFX2 U6911 ( .A(n2304), .Y(n6094) );
  AND2X1 U6912 ( .A(a_length[7]), .B(n8952), .Y(n3112) );
  INVX1 U6913 ( .A(n3112), .Y(n6095) );
  AND2X1 U6914 ( .A(a_length[18]), .B(n8953), .Y(n3090) );
  INVX1 U6915 ( .A(n3090), .Y(n6096) );
  AND2X1 U6916 ( .A(v_length[0]), .B(n8954), .Y(n2998) );
  INVX1 U6917 ( .A(n2998), .Y(n6097) );
  AND2X1 U6918 ( .A(v_length[9]), .B(n8955), .Y(n2980) );
  INVX1 U6919 ( .A(n2980), .Y(n6098) );
  AND2X1 U6920 ( .A(recentdatapoints_head_i[12]), .B(n8980), .Y(n1971) );
  INVX1 U6921 ( .A(n1971), .Y(n6099) );
  AND2X1 U6922 ( .A(recentdatapoints_head_i[20]), .B(n8979), .Y(n1963) );
  INVX1 U6923 ( .A(n1963), .Y(n6100) );
  AND2X1 U6924 ( .A(CircularBuffer_head_i_read_ass_reg_1624[6]), .B(n9011), 
        .Y(n1787) );
  INVX1 U6925 ( .A(n1787), .Y(n6101) );
  AND2X1 U6926 ( .A(CircularBuffer_head_i_read_ass_reg_1624[13]), .B(n9010), 
        .Y(n1766) );
  INVX1 U6927 ( .A(n1766), .Y(n6102) );
  AND2X1 U6928 ( .A(CircularBuffer_head_i_read_ass_reg_1624[20]), .B(n9009), 
        .Y(n1745) );
  INVX1 U6929 ( .A(n1745), .Y(n6103) );
  AND2X1 U6930 ( .A(n2794), .B(n8992), .Y(n1648) );
  INVX1 U6931 ( .A(n1648), .Y(n6104) );
  AND2X1 U6932 ( .A(n2782), .B(n8991), .Y(n1639) );
  INVX1 U6933 ( .A(n1639), .Y(n6105) );
  AND2X1 U6934 ( .A(n2762), .B(n8993), .Y(n1624) );
  INVX1 U6935 ( .A(n1624), .Y(n6106) );
  BUFX2 U6936 ( .A(n2857), .Y(n6107) );
  BUFX2 U6937 ( .A(n2833), .Y(n6108) );
  AND2X1 U6938 ( .A(CircularBuffer_sum_read_assign_reg_1610[7]), .B(n9006), 
        .Y(n1452) );
  INVX1 U6939 ( .A(n1452), .Y(n6109) );
  AND2X1 U6940 ( .A(n9012), .B(sum_phi_fu_311_p4[3]), .Y(n2684) );
  INVX1 U6941 ( .A(n2684), .Y(n6110) );
  BUFX2 U6942 ( .A(n2728), .Y(n6111) );
  AND2X1 U6943 ( .A(n9012), .B(sum_phi_fu_311_p4[17]), .Y(n2628) );
  INVX1 U6944 ( .A(n2628), .Y(n6112) );
  BUFX2 U6945 ( .A(n2715), .Y(n6113) );
  AND2X1 U6946 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[18]), .B(n9033), 
        .Y(n1376) );
  INVX1 U6947 ( .A(n1376), .Y(n6114) );
  AND2X1 U6948 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[8]), .B(n9035), 
        .Y(n1356) );
  INVX1 U6949 ( .A(n1356), .Y(n6115) );
  AND2X1 U6950 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[4]), .B(n9036), 
        .Y(n1348) );
  INVX1 U6951 ( .A(n1348), .Y(n6116) );
  AND2X1 U6952 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[8]), .B(n9038), 
        .Y(n1326) );
  INVX1 U6953 ( .A(n1326), .Y(n6117) );
  AND2X1 U6954 ( .A(recentABools_head_i[10]), .B(n9039), .Y(n1319) );
  INVX1 U6955 ( .A(n1319), .Y(n6118) );
  AND2X1 U6956 ( .A(recentABools_head_i[31]), .B(n9037), .Y(n1270) );
  INVX1 U6957 ( .A(n1270), .Y(n6119) );
  AND2X1 U6958 ( .A(VbeatFallDelay_new_1_reg_342[8]), .B(n9013), .Y(n2165) );
  INVX1 U6959 ( .A(n2165), .Y(n6120) );
  AND2X1 U6960 ( .A(tmp_5_fu_726_p2[22]), .B(n8994), .Y(n1120) );
  INVX1 U6961 ( .A(n1120), .Y(n6121) );
  AND2X1 U6962 ( .A(tmp_4_fu_716_p2[9]), .B(n8995), .Y(n1050) );
  INVX1 U6963 ( .A(n1050), .Y(n6122) );
  AND2X1 U6964 ( .A(tmp_4_fu_716_p2[28]), .B(n8996), .Y(n985) );
  INVX1 U6965 ( .A(n985), .Y(n6123) );
  AND2X1 U6966 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[1]), .Y(n2410) );
  INVX1 U6967 ( .A(n2410), .Y(n6124) );
  AND2X1 U6968 ( .A(AbeatDelay[8]), .B(n10670), .Y(n764) );
  INVX1 U6969 ( .A(n764), .Y(n6125) );
  AND2X1 U6970 ( .A(AbeatDelay_new_reg_394[11]), .B(n9041), .Y(n2223) );
  INVX1 U6971 ( .A(n2223), .Y(n6126) );
  AND2X1 U6972 ( .A(tmp_3_fu_706_p2[15]), .B(n8997), .Y(n743) );
  INVX1 U6973 ( .A(n743), .Y(n6127) );
  AND2X1 U6974 ( .A(AbeatDelay[21]), .B(n10670), .Y(n720) );
  INVX1 U6975 ( .A(n720), .Y(n6128) );
  AND2X1 U6976 ( .A(AstimDelay[8]), .B(n8896), .Y(n659) );
  INVX1 U6977 ( .A(n659), .Y(n6129) );
  AND2X1 U6978 ( .A(tmp_6_fu_497_p3[12]), .B(n8966), .Y(n648) );
  INVX1 U6979 ( .A(n648), .Y(n6130) );
  AND2X1 U6980 ( .A(AstimDelay[25]), .B(n8896), .Y(n608) );
  INVX1 U6981 ( .A(n608), .Y(n6131) );
  AND2X1 U6982 ( .A(VstimDelay[11]), .B(n10670), .Y(n550) );
  INVX1 U6983 ( .A(n550), .Y(n6132) );
  AND2X1 U6984 ( .A(tmp_7_fu_511_p3[14]), .B(n8964), .Y(n542) );
  INVX1 U6985 ( .A(n542), .Y(n6133) );
  AND2X1 U6986 ( .A(\Decision_AXILiteS_s_axi_U/n368 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n415 ) );
  INVX1 U6987 ( .A(\Decision_AXILiteS_s_axi_U/n415 ), .Y(n6134) );
  AND2X1 U6988 ( .A(\Decision_AXILiteS_s_axi_U/n564 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n521 ) );
  INVX1 U6989 ( .A(\Decision_AXILiteS_s_axi_U/n521 ), .Y(n6135) );
  AND2X1 U6990 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[3]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n385 )
         );
  INVX1 U6991 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n385 ), 
        .Y(n6136) );
  AND2X1 U6992 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[9]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n397 )
         );
  INVX1 U6993 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n397 ), 
        .Y(n6137) );
  AND2X1 U6994 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[6]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n426 )
         );
  INVX1 U6995 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n426 ), 
        .Y(n6138) );
  AND2X1 U6996 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[7]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n462 )
         );
  INVX1 U6997 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n462 ), 
        .Y(n6139) );
  AND2X1 U6998 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[0]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n482 )
         );
  INVX1 U6999 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n482 ), 
        .Y(n6140) );
  AND2X1 U7000 ( .A(n9467), .B(data_read_reg_1495[1]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n518 )
         );
  INVX1 U7001 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n518 ), 
        .Y(n6141) );
  AND2X1 U7002 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][11] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n573 )
         );
  INVX1 U7003 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n573 ), 
        .Y(n6142) );
  AND2X1 U7004 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][8] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n661 )
         );
  INVX1 U7005 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n661 ), 
        .Y(n6143) );
  AND2X1 U7006 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][9] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n681 )
         );
  INVX1 U7007 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n681 ), 
        .Y(n6144) );
  AND2X1 U7008 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][6] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n696 )
         );
  INVX1 U7009 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n696 ), 
        .Y(n6145) );
  AND2X1 U7010 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][7] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n714 )
         );
  INVX1 U7011 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n714 ), 
        .Y(n6146) );
  AND2X1 U7012 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][4] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n728 )
         );
  INVX1 U7013 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n728 ), 
        .Y(n6147) );
  AND2X1 U7014 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][5] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n746 )
         );
  INVX1 U7015 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n746 ), 
        .Y(n6148) );
  AND2X1 U7016 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][2] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n760 )
         );
  INVX1 U7017 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n760 ), 
        .Y(n6149) );
  AND2X1 U7018 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][3] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n812 )
         );
  INVX1 U7019 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n812 ), 
        .Y(n6150) );
  AND2X1 U7020 ( .A(sum_reg_308[23]), .B(n8929), .Y(n2606) );
  INVX1 U7021 ( .A(n2606), .Y(n6151) );
  AND2X1 U7022 ( .A(sum_1_reg_376[7]), .B(n8930), .Y(n2436) );
  INVX1 U7023 ( .A(n2436), .Y(n6152) );
  AND2X1 U7024 ( .A(tmp_29_i_fu_752_p2[24]), .B(n8920), .Y(n3168) );
  INVX1 U7025 ( .A(n3168), .Y(n6153) );
  AND2X1 U7026 ( .A(tmp_29_i1_fu_1065_p2[24]), .B(n8922), .Y(n3220) );
  INVX1 U7027 ( .A(n3220), .Y(n6154) );
  INVX1 U7028 ( .A(n4625), .Y(n6155) );
  AND2X1 U7029 ( .A(ACaptureThresh_loc_reg_288[9]), .B(n8970), .Y(n3044) );
  INVX1 U7030 ( .A(n3044), .Y(n6156) );
  BUFX2 U7031 ( .A(n3043), .Y(n6157) );
  INVX1 U7032 ( .A(n4615), .Y(n6158) );
  AND2X1 U7033 ( .A(ACaptureThresh_loc_reg_288[19]), .B(n8971), .Y(n3024) );
  INVX1 U7034 ( .A(n3024), .Y(n6159) );
  BUFX2 U7035 ( .A(n3023), .Y(n6160) );
  INVX1 U7036 ( .A(n4554), .Y(n6161) );
  AND2X1 U7037 ( .A(VCaptureThresh_loc_reg_298[16]), .B(n8969), .Y(n2902) );
  INVX1 U7038 ( .A(n2902), .Y(n6162) );
  BUFX2 U7039 ( .A(n2901), .Y(n6163) );
  AND2X1 U7040 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[7]), 
        .Y(n446) );
  INVX1 U7041 ( .A(n446), .Y(n6164) );
  AND2X1 U7042 ( .A(CircularBuffer_len_read_assign_fu_772_p2[29]), .B(n8919), 
        .Y(n2736) );
  INVX1 U7043 ( .A(n2736), .Y(n6165) );
  AND2X1 U7044 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[29]), .B(n8921), .Y(n2243) );
  INVX1 U7045 ( .A(n2243), .Y(n6166) );
  AND2X1 U7046 ( .A(v_flip[4]), .B(n8952), .Y(n3132) );
  INVX1 U7047 ( .A(n3132), .Y(n6167) );
  AND2X1 U7048 ( .A(a_length[19]), .B(n8953), .Y(n3088) );
  INVX1 U7049 ( .A(n3088), .Y(n6168) );
  AND2X1 U7050 ( .A(v_length[4]), .B(n8954), .Y(n2990) );
  INVX1 U7051 ( .A(n2990), .Y(n6169) );
  AND2X1 U7052 ( .A(v_length[10]), .B(n8955), .Y(n2978) );
  INVX1 U7053 ( .A(n2978), .Y(n6170) );
  AND2X1 U7054 ( .A(recentdatapoints_head_i[7]), .B(n8980), .Y(n1976) );
  INVX1 U7055 ( .A(n1976), .Y(n6171) );
  AND2X1 U7056 ( .A(recentdatapoints_head_i[21]), .B(n8979), .Y(n1962) );
  INVX1 U7057 ( .A(n1962), .Y(n6172) );
  AND2X1 U7058 ( .A(recentdatapoints_head_i[22]), .B(n8980), .Y(n1961) );
  INVX1 U7059 ( .A(n1961), .Y(n6173) );
  AND2X1 U7060 ( .A(recentVBools_head_i[6]), .B(n9011), .Y(n1786) );
  INVX1 U7061 ( .A(n1786), .Y(n6174) );
  AND2X1 U7062 ( .A(recentVBools_head_i[13]), .B(n9010), .Y(n1765) );
  INVX1 U7063 ( .A(n1765), .Y(n6175) );
  AND2X1 U7064 ( .A(recentVBools_head_i[20]), .B(n9009), .Y(n1744) );
  INVX1 U7065 ( .A(n1744), .Y(n6176) );
  BUFX2 U7066 ( .A(n2735), .Y(n6177) );
  AND2X1 U7067 ( .A(n2780), .B(n8992), .Y(n1638) );
  INVX1 U7068 ( .A(n1638), .Y(n6178) );
  AND2X1 U7069 ( .A(n2760), .B(n8993), .Y(n1623) );
  INVX1 U7070 ( .A(n1623), .Y(n6179) );
  BUFX2 U7071 ( .A(n2855), .Y(n6180) );
  BUFX2 U7072 ( .A(n2831), .Y(n6181) );
  AND2X1 U7073 ( .A(CircularBuffer_sum_read_assign_reg_1610[1]), .B(n9007), 
        .Y(n1464) );
  INVX1 U7074 ( .A(n1464), .Y(n6182) );
  AND2X1 U7075 ( .A(CircularBuffer_sum_read_assign_reg_1610[8]), .B(n9006), 
        .Y(n1450) );
  INVX1 U7076 ( .A(n1450), .Y(n6183) );
  AND2X1 U7077 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[4]), .Y(n2680) );
  INVX1 U7078 ( .A(n2680), .Y(n6184) );
  BUFX2 U7079 ( .A(n2727), .Y(n6185) );
  AND2X1 U7080 ( .A(n9012), .B(sum_phi_fu_311_p4[18]), .Y(n2624) );
  INVX1 U7081 ( .A(n2624), .Y(n6186) );
  BUFX2 U7082 ( .A(n2714), .Y(n6187) );
  AND2X1 U7083 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[3]), .B(n9036), 
        .Y(n1346) );
  INVX1 U7084 ( .A(n1346), .Y(n6188) );
  AND2X1 U7085 ( .A(n10271), .B(n9019), .Y(n1338) );
  INVX1 U7086 ( .A(n1338), .Y(n6189) );
  AND2X1 U7087 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[7]), .B(n9038), 
        .Y(n1328) );
  INVX1 U7088 ( .A(n1328), .Y(n6190) );
  AND2X1 U7089 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[10]), .B(n9039), 
        .Y(n1320) );
  INVX1 U7090 ( .A(n1320), .Y(n6191) );
  AND2X1 U7091 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[12]), .B(n9040), 
        .Y(n1315) );
  INVX1 U7092 ( .A(n1315), .Y(n6192) );
  AND2X1 U7093 ( .A(VbeatFallDelay[0]), .B(n9037), .Y(n1208) );
  INVX1 U7094 ( .A(n1208), .Y(n6193) );
  AND2X1 U7095 ( .A(VbeatFallDelay_new_1_reg_342[1]), .B(n9013), .Y(n2158) );
  INVX1 U7096 ( .A(n2158), .Y(n6194) );
  AND2X1 U7097 ( .A(VbeatFallDelay_new_1_reg_342[15]), .B(n9013), .Y(n2172) );
  INVX1 U7098 ( .A(n2172), .Y(n6195) );
  AND2X1 U7099 ( .A(tmp_5_fu_726_p2[23]), .B(n8994), .Y(n1116) );
  INVX1 U7100 ( .A(n1116), .Y(n6196) );
  AND2X1 U7101 ( .A(VbeatFallDelay[23]), .B(n9035), .Y(n1114) );
  INVX1 U7102 ( .A(n1114), .Y(n6197) );
  AND2X1 U7103 ( .A(tmp_4_fu_716_p2[10]), .B(n8995), .Y(n1047) );
  INVX1 U7104 ( .A(n1047), .Y(n6198) );
  AND2X1 U7105 ( .A(tmp_4_fu_716_p2[29]), .B(n8996), .Y(n981) );
  INVX1 U7106 ( .A(n981), .Y(n6199) );
  AND2X1 U7107 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[0]), .Y(n2406) );
  INVX1 U7108 ( .A(n2406), .Y(n6200) );
  BUFX2 U7109 ( .A(n2330), .Y(n6201) );
  AND2X1 U7110 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[8]), .Y(n2438) );
  INVX1 U7111 ( .A(n2438), .Y(n6202) );
  BUFX2 U7112 ( .A(n2317), .Y(n6203) );
  BUFX2 U7113 ( .A(n2374), .Y(n6204) );
  AND2X1 U7114 ( .A(AbeatDelay[10]), .B(n10670), .Y(n758) );
  INVX1 U7115 ( .A(n758), .Y(n6205) );
  AND2X1 U7116 ( .A(AbeatDelay_new_reg_394[12]), .B(n9041), .Y(n2222) );
  INVX1 U7117 ( .A(n2222), .Y(n6206) );
  AND2X1 U7118 ( .A(tmp_3_fu_706_p2[16]), .B(n8997), .Y(n739) );
  INVX1 U7119 ( .A(n739), .Y(n6207) );
  AND2X1 U7120 ( .A(AbeatDelay[25]), .B(n8896), .Y(n706) );
  INVX1 U7121 ( .A(n706), .Y(n6208) );
  AND2X1 U7122 ( .A(AstimDelay[9]), .B(n8896), .Y(n656) );
  INVX1 U7123 ( .A(n656), .Y(n6209) );
  AND2X1 U7124 ( .A(tmp_6_fu_497_p3[18]), .B(n8966), .Y(n630) );
  INVX1 U7125 ( .A(n630), .Y(n6210) );
  AND2X1 U7126 ( .A(AstimDelay[26]), .B(n10670), .Y(n605) );
  INVX1 U7127 ( .A(n605), .Y(n6211) );
  AND2X1 U7128 ( .A(VstimDelay[12]), .B(n10670), .Y(n547) );
  INVX1 U7129 ( .A(n547), .Y(n6212) );
  AND2X1 U7130 ( .A(tmp_7_fu_511_p3[15]), .B(n8964), .Y(n539) );
  INVX1 U7131 ( .A(n539), .Y(n6213) );
  AND2X1 U7132 ( .A(\Decision_AXILiteS_s_axi_U/n364 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n413 ) );
  INVX1 U7133 ( .A(\Decision_AXILiteS_s_axi_U/n413 ), .Y(n6214) );
  AND2X1 U7134 ( .A(\Decision_AXILiteS_s_axi_U/n366 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n456 ) );
  INVX1 U7135 ( .A(\Decision_AXILiteS_s_axi_U/n456 ), .Y(n6215) );
  AND2X1 U7136 ( .A(\Decision_AXILiteS_s_axi_U/n368 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n520 ) );
  INVX1 U7137 ( .A(\Decision_AXILiteS_s_axi_U/n520 ), .Y(n6216) );
  AND2X1 U7138 ( .A(\Decision_AXILiteS_s_axi_U/n564 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n563 ) );
  INVX1 U7139 ( .A(\Decision_AXILiteS_s_axi_U/n563 ), .Y(n6217) );
  AND2X1 U7140 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[4]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n387 )
         );
  INVX1 U7141 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n387 ), 
        .Y(n6218) );
  AND2X1 U7142 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[10]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n399 )
         );
  INVX1 U7143 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n399 ), 
        .Y(n6219) );
  AND2X1 U7144 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[1]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n416 )
         );
  INVX1 U7145 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n416 ), 
        .Y(n6220) );
  AND2X1 U7146 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[0]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n448 )
         );
  INVX1 U7147 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n448 ), 
        .Y(n6221) );
  AND2X1 U7148 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[7]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n496 )
         );
  INVX1 U7149 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n496 ), 
        .Y(n6222) );
  AND2X1 U7150 ( .A(n9467), .B(data_read_reg_1495[6]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n528 )
         );
  INVX1 U7151 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n528 ), 
        .Y(n6223) );
  AND2X1 U7152 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][8] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n567 )
         );
  INVX1 U7153 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n567 ), 
        .Y(n6224) );
  AND2X1 U7154 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][11] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n664 )
         );
  INVX1 U7155 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n664 ), 
        .Y(n6225) );
  AND2X1 U7156 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][10] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n682 )
         );
  INVX1 U7157 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n682 ), 
        .Y(n6226) );
  AND2X1 U7158 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][5] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n695 )
         );
  INVX1 U7159 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n695 ), 
        .Y(n6227) );
  AND2X1 U7160 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][4] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n711 )
         );
  INVX1 U7161 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n711 ), 
        .Y(n6228) );
  AND2X1 U7162 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][7] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n731 )
         );
  INVX1 U7163 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n731 ), 
        .Y(n6229) );
  AND2X1 U7164 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][6] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n747 )
         );
  INVX1 U7165 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n747 ), 
        .Y(n6230) );
  AND2X1 U7166 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][3] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n830 )
         );
  INVX1 U7167 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n830 ), 
        .Y(n6231) );
  AND2X1 U7168 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][2] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n846 )
         );
  INVX1 U7169 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n846 ), 
        .Y(n6232) );
  AND2X1 U7170 ( .A(tmp_29_i_fu_752_p2[30]), .B(n8920), .Y(n3161) );
  INVX1 U7171 ( .A(n3161), .Y(n6233) );
  AND2X1 U7172 ( .A(tmp_29_i1_fu_1065_p2[30]), .B(n8922), .Y(n3213) );
  INVX1 U7173 ( .A(n3213), .Y(n6234) );
  AND2X1 U7174 ( .A(sum_reg_308[0]), .B(n8929), .Y(n2698) );
  INVX1 U7175 ( .A(n2698), .Y(n6235) );
  AND2X1 U7176 ( .A(sum_reg_308[15]), .B(n8929), .Y(n2638) );
  INVX1 U7177 ( .A(n2638), .Y(n6236) );
  AND2X1 U7178 ( .A(sum_1_reg_376[27]), .B(n8930), .Y(n2516) );
  INVX1 U7179 ( .A(n2516), .Y(n6237) );
  AND2X1 U7180 ( .A(tmp_29_i_fu_752_p2[23]), .B(n8920), .Y(n3169) );
  INVX1 U7181 ( .A(n3169), .Y(n6238) );
  AND2X1 U7182 ( .A(tmp_29_i1_fu_1065_p2[23]), .B(n8922), .Y(n3221) );
  INVX1 U7183 ( .A(n3221), .Y(n6239) );
  INVX1 U7184 ( .A(n4630), .Y(n6240) );
  AND2X1 U7185 ( .A(ACaptureThresh_loc_reg_288[4]), .B(n8970), .Y(n3054) );
  INVX1 U7186 ( .A(n3054), .Y(n6241) );
  BUFX2 U7187 ( .A(n3053), .Y(n6242) );
  INVX1 U7188 ( .A(n4614), .Y(n6243) );
  AND2X1 U7189 ( .A(ACaptureThresh_loc_reg_288[20]), .B(n8971), .Y(n3022) );
  INVX1 U7190 ( .A(n3022), .Y(n6244) );
  BUFX2 U7191 ( .A(n3021), .Y(n6245) );
  INVX1 U7192 ( .A(n4568), .Y(n6246) );
  AND2X1 U7193 ( .A(VCaptureThresh_loc_reg_298[2]), .B(n8970), .Y(n2930) );
  INVX1 U7194 ( .A(n2930), .Y(n6247) );
  BUFX2 U7195 ( .A(n2929), .Y(n6248) );
  INVX1 U7196 ( .A(n4553), .Y(n6249) );
  AND2X1 U7197 ( .A(VCaptureThresh_loc_reg_298[17]), .B(n8969), .Y(n2900) );
  INVX1 U7198 ( .A(n2900), .Y(n6250) );
  BUFX2 U7199 ( .A(n2899), .Y(n6251) );
  AND2X1 U7200 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[14]), 
        .Y(n461) );
  INVX1 U7201 ( .A(n461), .Y(n6252) );
  AND2X1 U7202 ( .A(CircularBuffer_len_read_assign_fu_772_p2[16]), .B(n8919), 
        .Y(n2762) );
  INVX1 U7203 ( .A(n2762), .Y(n6253) );
  AND2X1 U7204 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[16]), .B(n8921), .Y(n2269) );
  INVX1 U7205 ( .A(n2269), .Y(n6254) );
  AND2X1 U7206 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[31]), .Y(n2530) );
  INVX1 U7207 ( .A(n2530), .Y(n6255) );
  AND2X1 U7208 ( .A(a_length[8]), .B(n8952), .Y(n3110) );
  INVX1 U7209 ( .A(n3110), .Y(n6256) );
  AND2X1 U7210 ( .A(a_length[20]), .B(n8953), .Y(n3086) );
  INVX1 U7211 ( .A(n3086), .Y(n6257) );
  AND2X1 U7212 ( .A(v_length[5]), .B(n8954), .Y(n2988) );
  INVX1 U7213 ( .A(n2988), .Y(n6258) );
  AND2X1 U7214 ( .A(v_length[11]), .B(n8955), .Y(n2976) );
  INVX1 U7215 ( .A(n2976), .Y(n6259) );
  AND2X1 U7216 ( .A(recentdatapoints_head_i[13]), .B(n8980), .Y(n1970) );
  INVX1 U7217 ( .A(n1970), .Y(n6260) );
  AND2X1 U7218 ( .A(recentdatapoints_head_i[29]), .B(n8979), .Y(n1954) );
  INVX1 U7219 ( .A(n1954), .Y(n6261) );
  AND2X1 U7220 ( .A(CircularBuffer_head_i_read_ass_reg_1624[7]), .B(n9011), 
        .Y(n1784) );
  INVX1 U7221 ( .A(n1784), .Y(n6262) );
  AND2X1 U7222 ( .A(CircularBuffer_head_i_read_ass_reg_1624[14]), .B(n9010), 
        .Y(n1763) );
  INVX1 U7223 ( .A(n1763), .Y(n6263) );
  AND2X1 U7224 ( .A(CircularBuffer_head_i_read_ass_reg_1624[21]), .B(n9009), 
        .Y(n1742) );
  INVX1 U7225 ( .A(n1742), .Y(n6264) );
  AND2X1 U7226 ( .A(recentVBools_head_i[29]), .B(n9008), .Y(n1717) );
  INVX1 U7227 ( .A(n1717), .Y(n6265) );
  AND2X1 U7228 ( .A(n2778), .B(n8992), .Y(n1637) );
  INVX1 U7229 ( .A(n1637), .Y(n6266) );
  BUFX2 U7230 ( .A(n2793), .Y(n6267) );
  BUFX2 U7231 ( .A(n2853), .Y(n6268) );
  BUFX2 U7232 ( .A(n2771), .Y(n6269) );
  BUFX2 U7233 ( .A(n2829), .Y(n6270) );
  AND2X1 U7234 ( .A(CircularBuffer_sum_read_assign_reg_1610[2]), .B(n9007), 
        .Y(n1462) );
  INVX1 U7235 ( .A(n1462), .Y(n6271) );
  AND2X1 U7236 ( .A(CircularBuffer_sum_read_assign_reg_1610[9]), .B(n9006), 
        .Y(n1448) );
  INVX1 U7237 ( .A(n1448), .Y(n6272) );
  AND2X1 U7238 ( .A(n9012), .B(sum_phi_fu_311_p4[5]), .Y(n2676) );
  INVX1 U7239 ( .A(n2676), .Y(n6273) );
  BUFX2 U7240 ( .A(n2726), .Y(n6274) );
  AND2X1 U7241 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[19]), .Y(n2620) );
  INVX1 U7242 ( .A(n2620), .Y(n6275) );
  BUFX2 U7243 ( .A(n2712), .Y(n6276) );
  AND2X1 U7244 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[26]), .B(n9032), 
        .Y(n1392) );
  INVX1 U7245 ( .A(n1392), .Y(n6277) );
  AND2X1 U7246 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[2]), .B(n9036), 
        .Y(n1344) );
  INVX1 U7247 ( .A(n1344), .Y(n6278) );
  AND2X1 U7248 ( .A(recentABools_head_i[7]), .B(n9038), .Y(n1327) );
  INVX1 U7249 ( .A(n1327), .Y(n6279) );
  AND2X1 U7250 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[11]), .B(n9039), 
        .Y(n1317) );
  INVX1 U7251 ( .A(n1317), .Y(n6280) );
  AND2X1 U7252 ( .A(recentABools_head_i[13]), .B(n9040), .Y(n1312) );
  INVX1 U7253 ( .A(n1312), .Y(n6281) );
  AND2X1 U7254 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[14]), .B(n9035), 
        .Y(n1311) );
  INVX1 U7255 ( .A(n1311), .Y(n6282) );
  AND2X1 U7256 ( .A(VbeatFallDelay[1]), .B(n9037), .Y(n1202) );
  INVX1 U7257 ( .A(n1202), .Y(n6283) );
  AND2X1 U7258 ( .A(VbeatFallDelay_new_1_reg_342[2]), .B(n9013), .Y(n2159) );
  INVX1 U7259 ( .A(n2159), .Y(n6284) );
  AND2X1 U7260 ( .A(tmp_5_fu_726_p2[6]), .B(n8993), .Y(n1184) );
  INVX1 U7261 ( .A(n1184), .Y(n6285) );
  AND2X1 U7262 ( .A(VbeatFallDelay_new_1_reg_342[16]), .B(n9013), .Y(n2173) );
  INVX1 U7263 ( .A(n2173), .Y(n6286) );
  AND2X1 U7264 ( .A(tmp_5_fu_726_p2[24]), .B(n8994), .Y(n1112) );
  INVX1 U7265 ( .A(n1112), .Y(n6287) );
  AND2X1 U7266 ( .A(VbeatFallDelay[25]), .B(n9034), .Y(n1106) );
  INVX1 U7267 ( .A(n1106), .Y(n6288) );
  AND2X1 U7268 ( .A(tmp_4_fu_716_p2[11]), .B(n8995), .Y(n1043) );
  INVX1 U7269 ( .A(n1043), .Y(n6289) );
  AND2X1 U7270 ( .A(tmp_4_fu_716_p2[30]), .B(n8996), .Y(n978) );
  INVX1 U7271 ( .A(n978), .Y(n6290) );
  AND2X1 U7272 ( .A(n2301), .B(n9019), .Y(n972) );
  INVX1 U7273 ( .A(n972), .Y(n6291) );
  AND2X1 U7274 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[9]), .Y(n2442) );
  INVX1 U7275 ( .A(n2442), .Y(n6292) );
  BUFX2 U7276 ( .A(n2322), .Y(n6293) );
  BUFX2 U7277 ( .A(n2316), .Y(n6294) );
  BUFX2 U7278 ( .A(n2398), .Y(n6295) );
  BUFX2 U7279 ( .A(n2298), .Y(n6296) );
  BUFX2 U7280 ( .A(n2370), .Y(n6297) );
  AND2X1 U7281 ( .A(AbeatDelay_new_reg_394[13]), .B(n9041), .Y(n2221) );
  INVX1 U7282 ( .A(n2221), .Y(n6298) );
  AND2X1 U7283 ( .A(AbeatDelay[13]), .B(n8896), .Y(n747) );
  INVX1 U7284 ( .A(n747), .Y(n6299) );
  AND2X1 U7285 ( .A(tmp_3_fu_706_p2[17]), .B(n8997), .Y(n735) );
  INVX1 U7286 ( .A(n735), .Y(n6300) );
  AND2X1 U7287 ( .A(AbeatDelay[26]), .B(n8896), .Y(n703) );
  INVX1 U7288 ( .A(n703), .Y(n6301) );
  AND2X1 U7289 ( .A(tmp_6_fu_497_p3[5]), .B(n8965), .Y(n669) );
  INVX1 U7290 ( .A(n669), .Y(n6302) );
  AND2X1 U7291 ( .A(AstimDelay[10]), .B(n8896), .Y(n653) );
  INVX1 U7292 ( .A(n653), .Y(n6303) );
  AND2X1 U7293 ( .A(tmp_6_fu_497_p3[19]), .B(n8966), .Y(n627) );
  INVX1 U7294 ( .A(n627), .Y(n6304) );
  AND2X1 U7295 ( .A(AstimDelay[27]), .B(n8896), .Y(n602) );
  INVX1 U7296 ( .A(n602), .Y(n6305) );
  AND2X1 U7297 ( .A(VstimDelay[13]), .B(n10670), .Y(n544) );
  INVX1 U7298 ( .A(n544), .Y(n6306) );
  AND2X1 U7299 ( .A(tmp_7_fu_511_p3[16]), .B(n8964), .Y(n536) );
  INVX1 U7300 ( .A(n536), .Y(n6307) );
  AND2X1 U7301 ( .A(\Decision_AXILiteS_s_axi_U/n362 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n412 ) );
  INVX1 U7302 ( .A(\Decision_AXILiteS_s_axi_U/n412 ), .Y(n6308) );
  AND2X1 U7303 ( .A(\Decision_AXILiteS_s_axi_U/n564 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n458 ) );
  INVX1 U7304 ( .A(\Decision_AXILiteS_s_axi_U/n458 ), .Y(n6309) );
  AND2X1 U7305 ( .A(\Decision_AXILiteS_s_axi_U/n366 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n519 ) );
  INVX1 U7306 ( .A(\Decision_AXILiteS_s_axi_U/n519 ), .Y(n6310) );
  AND2X1 U7307 ( .A(\Decision_AXILiteS_s_axi_U/n368 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n562 ) );
  INVX1 U7308 ( .A(\Decision_AXILiteS_s_axi_U/n562 ), .Y(n6311) );
  AND2X1 U7309 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[5]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n389 )
         );
  INVX1 U7310 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n389 ), 
        .Y(n6312) );
  AND2X1 U7311 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[11]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n401 )
         );
  INVX1 U7312 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n401 ), 
        .Y(n6313) );
  AND2X1 U7313 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[0]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n414 )
         );
  INVX1 U7314 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n414 ), 
        .Y(n6314) );
  AND2X1 U7315 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[1]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n450 )
         );
  INVX1 U7316 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n450 ), 
        .Y(n6315) );
  AND2X1 U7317 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[6]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n494 )
         );
  INVX1 U7318 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n494 ), 
        .Y(n6316) );
  AND2X1 U7319 ( .A(n9467), .B(data_read_reg_1495[7]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n530 )
         );
  INVX1 U7320 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n530 ), 
        .Y(n6317) );
  AND2X1 U7321 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][9] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n569 )
         );
  INVX1 U7322 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n569 ), 
        .Y(n6318) );
  AND2X1 U7323 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][10] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n663 )
         );
  INVX1 U7324 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n663 ), 
        .Y(n6319) );
  AND2X1 U7325 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][11] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n683 )
         );
  INVX1 U7326 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n683 ), 
        .Y(n6320) );
  AND2X1 U7327 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][4] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n694 )
         );
  INVX1 U7328 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n694 ), 
        .Y(n6321) );
  AND2X1 U7329 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][5] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n712 )
         );
  INVX1 U7330 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n712 ), 
        .Y(n6322) );
  AND2X1 U7331 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][6] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n730 )
         );
  INVX1 U7332 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n730 ), 
        .Y(n6323) );
  AND2X1 U7333 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][7] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n748 )
         );
  INVX1 U7334 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n748 ), 
        .Y(n6324) );
  AND2X1 U7335 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][2] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n829 )
         );
  INVX1 U7336 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n829 ), 
        .Y(n6325) );
  AND2X1 U7337 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][3] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n847 )
         );
  INVX1 U7338 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n847 ), 
        .Y(n6326) );
  AND2X1 U7339 ( .A(sum_1_reg_376[28]), .B(n8930), .Y(n2520) );
  INVX1 U7340 ( .A(n2520), .Y(n6327) );
  AND2X1 U7341 ( .A(sum_reg_308[2]), .B(n8929), .Y(n2690) );
  INVX1 U7342 ( .A(n2690), .Y(n6328) );
  AND2X1 U7343 ( .A(sum_reg_308[20]), .B(n8929), .Y(n2618) );
  INVX1 U7344 ( .A(n2618), .Y(n6329) );
  AND2X1 U7345 ( .A(sum_1_reg_376[24]), .B(n8930), .Y(n2504) );
  INVX1 U7346 ( .A(n2504), .Y(n6330) );
  AND2X1 U7347 ( .A(tmp_29_i_fu_752_p2[22]), .B(n8920), .Y(n3170) );
  INVX1 U7348 ( .A(n3170), .Y(n6331) );
  AND2X1 U7349 ( .A(tmp_29_i1_fu_1065_p2[22]), .B(n8922), .Y(n3222) );
  INVX1 U7350 ( .A(n3222), .Y(n6332) );
  AND2X1 U7351 ( .A(tmp_29_i_fu_752_p2[17]), .B(n8920), .Y(n3176) );
  INVX1 U7352 ( .A(n3176), .Y(n6333) );
  AND2X1 U7353 ( .A(tmp_29_i1_fu_1065_p2[17]), .B(n8922), .Y(n3228) );
  INVX1 U7354 ( .A(n3228), .Y(n6334) );
  INVX1 U7355 ( .A(n4629), .Y(n6335) );
  AND2X1 U7356 ( .A(ACaptureThresh_loc_reg_288[5]), .B(n8969), .Y(n3052) );
  INVX1 U7357 ( .A(n3052), .Y(n6336) );
  BUFX2 U7358 ( .A(n3051), .Y(n6337) );
  INVX1 U7359 ( .A(n4613), .Y(n6338) );
  AND2X1 U7360 ( .A(ACaptureThresh_loc_reg_288[21]), .B(n8971), .Y(n3020) );
  INVX1 U7361 ( .A(n3020), .Y(n6339) );
  BUFX2 U7362 ( .A(n3019), .Y(n6340) );
  INVX1 U7363 ( .A(n4567), .Y(n6341) );
  AND2X1 U7364 ( .A(VCaptureThresh_loc_reg_298[3]), .B(n8970), .Y(n2928) );
  INVX1 U7365 ( .A(n2928), .Y(n6342) );
  BUFX2 U7366 ( .A(n2927), .Y(n6343) );
  INVX1 U7367 ( .A(n4552), .Y(n6344) );
  AND2X1 U7368 ( .A(VCaptureThresh_loc_reg_298[18]), .B(n8969), .Y(n2898) );
  INVX1 U7369 ( .A(n2898), .Y(n6345) );
  BUFX2 U7370 ( .A(n2897), .Y(n6346) );
  AND2X1 U7371 ( .A(n9825), .B(n8972), .Y(n1988) );
  INVX1 U7372 ( .A(n1988), .Y(n6347) );
  AND2X1 U7373 ( .A(recentdatapoints_len_load_op_fu_556_p2[15]), .B(n8972), 
        .Y(n1837) );
  INVX1 U7374 ( .A(n1837), .Y(n6348) );
  AND2X1 U7375 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[10]), 
        .Y(n469) );
  INVX1 U7376 ( .A(n469), .Y(n6349) );
  AND2X1 U7377 ( .A(CircularBuffer_len_read_assign_fu_772_p2[17]), .B(n8919), 
        .Y(n2760) );
  INVX1 U7378 ( .A(n2760), .Y(n6350) );
  AND2X1 U7379 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[17]), .B(n8921), .Y(n2267) );
  INVX1 U7380 ( .A(n2267), .Y(n6351) );
  AND2X1 U7381 ( .A(a_flip[5]), .B(n8951), .Y(n3142) );
  INVX1 U7382 ( .A(n3142), .Y(n6352) );
  AND2X1 U7383 ( .A(a_length[21]), .B(n8953), .Y(n3084) );
  INVX1 U7384 ( .A(n3084), .Y(n6353) );
  AND2X1 U7385 ( .A(v_length[2]), .B(n8954), .Y(n2994) );
  INVX1 U7386 ( .A(n2994), .Y(n6354) );
  AND2X1 U7387 ( .A(v_length[12]), .B(n8955), .Y(n2974) );
  INVX1 U7388 ( .A(n2974), .Y(n6355) );
  AND2X1 U7389 ( .A(n8963), .B(recentdatapoints_head_i[3]), .Y(n1980) );
  INVX1 U7390 ( .A(n1980), .Y(n6356) );
  AND2X1 U7391 ( .A(recentdatapoints_head_i[10]), .B(n8977), .Y(n1973) );
  INVX1 U7392 ( .A(n1973), .Y(n6357) );
  AND2X1 U7393 ( .A(p_tmp_i_reg_1556[29]), .B(n8979), .Y(n1920) );
  INVX1 U7394 ( .A(n1920), .Y(n6358) );
  AND2X1 U7395 ( .A(p_tmp_i_reg_1556[17]), .B(n8980), .Y(n1896) );
  INVX1 U7396 ( .A(n1896), .Y(n6359) );
  AND2X1 U7397 ( .A(recentVBools_head_i[7]), .B(n9011), .Y(n1783) );
  INVX1 U7398 ( .A(n1783), .Y(n6360) );
  AND2X1 U7399 ( .A(recentVBools_head_i[15]), .B(n9010), .Y(n1759) );
  INVX1 U7400 ( .A(n1759), .Y(n6361) );
  AND2X1 U7401 ( .A(recentVBools_head_i[21]), .B(n9009), .Y(n1741) );
  INVX1 U7402 ( .A(n1741), .Y(n6362) );
  AND2X1 U7403 ( .A(CircularBuffer_head_i_read_ass_reg_1624[30]), .B(n9008), 
        .Y(n1715) );
  INVX1 U7404 ( .A(n1715), .Y(n6363) );
  BUFX2 U7405 ( .A(n2801), .Y(n6364) );
  AND2X1 U7406 ( .A(n2758), .B(n8992), .Y(n1622) );
  INVX1 U7407 ( .A(n1622), .Y(n6365) );
  AND2X1 U7408 ( .A(n2744), .B(n8991), .Y(n1612) );
  INVX1 U7409 ( .A(n1612), .Y(n6366) );
  BUFX2 U7410 ( .A(n2791), .Y(n6367) );
  BUFX2 U7411 ( .A(n2851), .Y(n6368) );
  BUFX2 U7412 ( .A(n2827), .Y(n6369) );
  BUFX2 U7413 ( .A(n2747), .Y(n6370) );
  AND2X1 U7414 ( .A(n8391), .B(n1646), .Y(n1602) );
  INVX1 U7415 ( .A(n1602), .Y(n6371) );
  AND2X1 U7416 ( .A(CircularBuffer_sum_read_assign_reg_1610[3]), .B(n9007), 
        .Y(n1460) );
  INVX1 U7417 ( .A(n1460), .Y(n6372) );
  AND2X1 U7418 ( .A(CircularBuffer_sum_read_assign_reg_1610[10]), .B(n9006), 
        .Y(n1446) );
  INVX1 U7419 ( .A(n1446), .Y(n6373) );
  AND2X1 U7420 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[6]), .Y(n2672) );
  INVX1 U7421 ( .A(n2672), .Y(n6374) );
  BUFX2 U7422 ( .A(n2725), .Y(n6375) );
  BUFX2 U7423 ( .A(n2713), .Y(n6376) );
  AND2X1 U7424 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[20]), .Y(n2616) );
  INVX1 U7425 ( .A(n2616), .Y(n6377) );
  AND2X1 U7426 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[20]), .B(n9032), 
        .Y(n1380) );
  INVX1 U7427 ( .A(n1380), .Y(n6378) );
  AND2X1 U7428 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[7]), .B(n9035), 
        .Y(n1354) );
  INVX1 U7429 ( .A(n1354), .Y(n6379) );
  AND2X1 U7430 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[1]), .B(n9036), 
        .Y(n1342) );
  INVX1 U7431 ( .A(n1342), .Y(n6380) );
  AND2X1 U7432 ( .A(recentABools_head_i[14]), .B(n9040), .Y(n1310) );
  INVX1 U7433 ( .A(n1310), .Y(n6381) );
  AND2X1 U7434 ( .A(recentABools_head_i[19]), .B(n9039), .Y(n1300) );
  INVX1 U7435 ( .A(n1300), .Y(n6382) );
  AND2X1 U7436 ( .A(recentABools_head_i[25]), .B(n9038), .Y(n1284) );
  INVX1 U7437 ( .A(n1284), .Y(n6383) );
  AND2X1 U7438 ( .A(VbeatFallDelay[2]), .B(n9037), .Y(n1198) );
  INVX1 U7439 ( .A(n1198), .Y(n6384) );
  AND2X1 U7440 ( .A(VbeatFallDelay_new_1_reg_342[3]), .B(n9013), .Y(n2160) );
  INVX1 U7441 ( .A(n2160), .Y(n6385) );
  AND2X1 U7442 ( .A(tmp_5_fu_726_p2[7]), .B(n8993), .Y(n1180) );
  INVX1 U7443 ( .A(n1180), .Y(n6386) );
  AND2X1 U7444 ( .A(VbeatFallDelay_new_1_reg_342[17]), .B(n9013), .Y(n2174) );
  INVX1 U7445 ( .A(n2174), .Y(n6387) );
  AND2X1 U7446 ( .A(tmp_5_fu_726_p2[25]), .B(n8994), .Y(n1108) );
  INVX1 U7447 ( .A(n1108), .Y(n6388) );
  AND2X1 U7448 ( .A(VbeatFallDelay[26]), .B(n9034), .Y(n1102) );
  INVX1 U7449 ( .A(n1102), .Y(n6389) );
  AND2X1 U7450 ( .A(VbeatDelay[1]), .B(n9033), .Y(n1073) );
  INVX1 U7451 ( .A(n1073), .Y(n6390) );
  AND2X1 U7452 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[8]), .Y(n2558) );
  INVX1 U7453 ( .A(n2558), .Y(n6391) );
  AND2X1 U7454 ( .A(tmp_4_fu_716_p2[12]), .B(n8995), .Y(n1039) );
  INVX1 U7455 ( .A(n1039), .Y(n6392) );
  AND2X1 U7456 ( .A(VbeatDelay[14]), .B(n9031), .Y(n1031) );
  INVX1 U7457 ( .A(n1031), .Y(n6393) );
  AND2X1 U7458 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[20]), .Y(n2546) );
  INVX1 U7459 ( .A(n2546), .Y(n6394) );
  AND2X1 U7460 ( .A(tmp_4_fu_716_p2[31]), .B(n8996), .Y(n975) );
  INVX1 U7461 ( .A(n975), .Y(n6395) );
  BUFX2 U7462 ( .A(n2329), .Y(n6396) );
  AND2X1 U7463 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[11]), .Y(n2450) );
  INVX1 U7464 ( .A(n2450), .Y(n6397) );
  BUFX2 U7465 ( .A(n2315), .Y(n6398) );
  AND2X1 U7466 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[22]), .Y(n2494) );
  INVX1 U7467 ( .A(n2494), .Y(n6399) );
  AND2X1 U7468 ( .A(n2287), .B(n9019), .Y(n962) );
  INVX1 U7469 ( .A(n962), .Y(n6400) );
  BUFX2 U7470 ( .A(n2396), .Y(n6401) );
  BUFX2 U7471 ( .A(n2292), .Y(n6402) );
  BUFX2 U7472 ( .A(n2368), .Y(n6403) );
  AND2X1 U7473 ( .A(n8392), .B(n970), .Y(n926) );
  INVX1 U7474 ( .A(n926), .Y(n6404) );
  AND2X1 U7475 ( .A(AbeatDelay[14]), .B(n8896), .Y(n744) );
  INVX1 U7476 ( .A(n744), .Y(n6405) );
  AND2X1 U7477 ( .A(tmp_3_fu_706_p2[18]), .B(n8997), .Y(n732) );
  INVX1 U7478 ( .A(n732), .Y(n6406) );
  AND2X1 U7479 ( .A(AbeatDelay_new_reg_394[19]), .B(n9041), .Y(n2215) );
  INVX1 U7480 ( .A(n2215), .Y(n6407) );
  AND2X1 U7481 ( .A(AbeatDelay[27]), .B(n10670), .Y(n700) );
  INVX1 U7482 ( .A(n700), .Y(n6408) );
  AND2X1 U7483 ( .A(AstimDelay[11]), .B(n8896), .Y(n650) );
  INVX1 U7484 ( .A(n650), .Y(n6409) );
  AND2X1 U7485 ( .A(tmp_6_fu_497_p3[13]), .B(n8966), .Y(n645) );
  INVX1 U7486 ( .A(n645), .Y(n6410) );
  AND2X1 U7487 ( .A(AstimDelay[28]), .B(n10670), .Y(n599) );
  INVX1 U7488 ( .A(n599), .Y(n6411) );
  AND2X1 U7489 ( .A(tmp_7_fu_511_p3[1]), .B(n8965), .Y(n581) );
  INVX1 U7490 ( .A(n581), .Y(n6412) );
  AND2X1 U7491 ( .A(VstimDelay[14]), .B(n10670), .Y(n541) );
  INVX1 U7492 ( .A(n541), .Y(n6413) );
  AND2X1 U7493 ( .A(tmp_7_fu_511_p3[17]), .B(n8964), .Y(n533) );
  INVX1 U7494 ( .A(n533), .Y(n6414) );
  AND2X1 U7495 ( .A(\Decision_AXILiteS_s_axi_U/n360 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n411 ) );
  INVX1 U7496 ( .A(\Decision_AXILiteS_s_axi_U/n411 ), .Y(n6415) );
  AND2X1 U7497 ( .A(\Decision_AXILiteS_s_axi_U/n368 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n457 ) );
  INVX1 U7498 ( .A(\Decision_AXILiteS_s_axi_U/n457 ), .Y(n6416) );
  AND2X1 U7499 ( .A(a_length[24]), .B(n8116), .Y(
        \Decision_AXILiteS_s_axi_U/n428 ) );
  INVX1 U7500 ( .A(\Decision_AXILiteS_s_axi_U/n428 ), .Y(n6417) );
  AND2X1 U7501 ( .A(\Decision_AXILiteS_s_axi_U/n364 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n518 ) );
  INVX1 U7502 ( .A(\Decision_AXILiteS_s_axi_U/n518 ), .Y(n6418) );
  AND2X1 U7503 ( .A(\Decision_AXILiteS_s_axi_U/n366 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n561 ) );
  INVX1 U7504 ( .A(\Decision_AXILiteS_s_axi_U/n561 ), .Y(n6419) );
  AND2X1 U7505 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[12]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n403 )
         );
  INVX1 U7506 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n403 ), 
        .Y(n6420) );
  AND2X1 U7507 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][14] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n579 )
         );
  INVX1 U7508 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n579 ), 
        .Y(n6421) );
  AND2X1 U7509 ( .A(n9468), .B(data_read_reg_1495[7]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n598 )
         );
  INVX1 U7510 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n598 ), 
        .Y(n6422) );
  AND2X1 U7511 ( .A(n9469), .B(data_read_reg_1495[6]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n630 )
         );
  INVX1 U7512 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n630 ), 
        .Y(n6423) );
  AND2X1 U7513 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][1] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n654 )
         );
  INVX1 U7514 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n654 ), 
        .Y(n6424) );
  AND2X1 U7515 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][13] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n666 )
         );
  INVX1 U7516 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n666 ), 
        .Y(n6425) );
  AND2X1 U7517 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][0] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n672 )
         );
  INVX1 U7518 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n672 ), 
        .Y(n6426) );
  AND2X1 U7519 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][12] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n684 )
         );
  INVX1 U7520 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n684 ), 
        .Y(n6427) );
  AND2X1 U7521 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][3] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n693 )
         );
  INVX1 U7522 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n693 ), 
        .Y(n6428) );
  AND2X1 U7523 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][2] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n709 )
         );
  INVX1 U7524 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n709 ), 
        .Y(n6429) );
  AND2X1 U7525 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][7] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n765 )
         );
  INVX1 U7526 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n765 ), 
        .Y(n6430) );
  AND2X1 U7527 ( .A(n9466), .B(data_read_reg_1495[1]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n778 )
         );
  INVX1 U7528 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n778 ), 
        .Y(n6431) );
  AND2X1 U7529 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][6] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n815 )
         );
  INVX1 U7530 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n815 ), 
        .Y(n6432) );
  AND2X1 U7531 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][5] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n832 )
         );
  INVX1 U7532 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n832 ), 
        .Y(n6433) );
  AND2X1 U7533 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][4] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n848 )
         );
  INVX1 U7534 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n848 ), 
        .Y(n6434) );
  AND2X1 U7535 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[0]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n862 )
         );
  INVX1 U7536 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n862 ), 
        .Y(n6435) );
  AND2X1 U7537 ( .A(sum_reg_308[11]), .B(n8929), .Y(n2654) );
  INVX1 U7538 ( .A(n2654), .Y(n6436) );
  AND2X1 U7539 ( .A(sum_1_reg_376[15]), .B(n8930), .Y(n2468) );
  INVX1 U7540 ( .A(n2468), .Y(n6437) );
  AND2X1 U7541 ( .A(sum_reg_308[24]), .B(n8929), .Y(n2602) );
  INVX1 U7542 ( .A(n2602), .Y(n6438) );
  AND2X1 U7543 ( .A(sum_1_reg_376[12]), .B(n8930), .Y(n2456) );
  INVX1 U7544 ( .A(n2456), .Y(n6439) );
  AND2X1 U7545 ( .A(tmp_29_i_fu_752_p2[21]), .B(n8920), .Y(n3171) );
  INVX1 U7546 ( .A(n3171), .Y(n6440) );
  AND2X1 U7547 ( .A(tmp_29_i1_fu_1065_p2[21]), .B(n8922), .Y(n3223) );
  INVX1 U7548 ( .A(n3223), .Y(n6441) );
  AND2X1 U7549 ( .A(tmp_29_i_fu_752_p2[12]), .B(n8920), .Y(n3181) );
  INVX1 U7550 ( .A(n3181), .Y(n6442) );
  AND2X1 U7551 ( .A(tmp_29_i1_fu_1065_p2[12]), .B(n8922), .Y(n3233) );
  INVX1 U7552 ( .A(n3233), .Y(n6443) );
  INVX1 U7553 ( .A(n4628), .Y(n6444) );
  AND2X1 U7554 ( .A(ACaptureThresh_loc_reg_288[6]), .B(n8970), .Y(n3050) );
  INVX1 U7555 ( .A(n3050), .Y(n6445) );
  BUFX2 U7556 ( .A(n3049), .Y(n6446) );
  INVX1 U7557 ( .A(n4612), .Y(n6447) );
  AND2X1 U7558 ( .A(ACaptureThresh_loc_reg_288[22]), .B(n8971), .Y(n3018) );
  INVX1 U7559 ( .A(n3018), .Y(n6448) );
  BUFX2 U7560 ( .A(n3017), .Y(n6449) );
  INVX1 U7561 ( .A(n4566), .Y(n6450) );
  AND2X1 U7562 ( .A(VCaptureThresh_loc_reg_298[4]), .B(n8970), .Y(n2926) );
  INVX1 U7563 ( .A(n2926), .Y(n6451) );
  BUFX2 U7564 ( .A(n2925), .Y(n6452) );
  INVX1 U7565 ( .A(n4550), .Y(n6453) );
  AND2X1 U7566 ( .A(VCaptureThresh_loc_reg_298[20]), .B(n8969), .Y(n2894) );
  INVX1 U7567 ( .A(n2894), .Y(n6454) );
  BUFX2 U7568 ( .A(n2893), .Y(n6455) );
  AND2X1 U7569 ( .A(recentdatapoints_len_load_op_fu_556_p2[10]), .B(n8972), 
        .Y(n1831) );
  INVX1 U7570 ( .A(n1831), .Y(n6456) );
  AND2X1 U7571 ( .A(recentdatapoints_len_load_op_fu_556_p2[16]), .B(n8972), 
        .Y(n1838) );
  INVX1 U7572 ( .A(n1838), .Y(n6457) );
  AND2X1 U7573 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[2]), 
        .Y(n456) );
  INVX1 U7574 ( .A(n456), .Y(n6458) );
  AND2X1 U7575 ( .A(CircularBuffer_len_read_assign_fu_772_p2[20]), .B(n8919), 
        .Y(n2754) );
  INVX1 U7576 ( .A(n2754), .Y(n6459) );
  AND2X1 U7577 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[20]), .B(n8921), .Y(n2261) );
  INVX1 U7578 ( .A(n2261), .Y(n6460) );
  AND2X1 U7579 ( .A(a_length[22]), .B(n8953), .Y(n3082) );
  INVX1 U7580 ( .A(n3082), .Y(n6461) );
  AND2X1 U7581 ( .A(v_length[3]), .B(n8954), .Y(n2992) );
  INVX1 U7582 ( .A(n2992), .Y(n6462) );
  AND2X1 U7583 ( .A(v_length[13]), .B(n8955), .Y(n2972) );
  INVX1 U7584 ( .A(n2972), .Y(n6463) );
  AND2X1 U7585 ( .A(v_length[14]), .B(n8952), .Y(n2970) );
  INVX1 U7586 ( .A(n2970), .Y(n6464) );
  AND2X1 U7587 ( .A(recentdatapoints_head_i[5]), .B(n8977), .Y(n1978) );
  INVX1 U7588 ( .A(n1978), .Y(n6465) );
  AND2X1 U7589 ( .A(recentdatapoints_head_i[23]), .B(n8978), .Y(n1960) );
  INVX1 U7590 ( .A(n1960), .Y(n6466) );
  AND2X1 U7591 ( .A(n8963), .B(recentdatapoints_head_i[2]), .Y(n1926) );
  INVX1 U7592 ( .A(n1926), .Y(n6467) );
  AND2X1 U7593 ( .A(p_tmp_i_reg_1556[28]), .B(n8979), .Y(n1918) );
  INVX1 U7594 ( .A(n1918), .Y(n6468) );
  AND2X1 U7595 ( .A(p_tmp_i_reg_1556[16]), .B(n8980), .Y(n1894) );
  INVX1 U7596 ( .A(n1894), .Y(n6469) );
  AND2X1 U7597 ( .A(CircularBuffer_head_i_read_ass_reg_1624[8]), .B(n9011), 
        .Y(n1781) );
  INVX1 U7598 ( .A(n1781), .Y(n6470) );
  AND2X1 U7599 ( .A(CircularBuffer_head_i_read_ass_reg_1624[16]), .B(n9010), 
        .Y(n1757) );
  INVX1 U7600 ( .A(n1757), .Y(n6471) );
  AND2X1 U7601 ( .A(CircularBuffer_head_i_read_ass_reg_1624[23]), .B(n9009), 
        .Y(n1736) );
  INVX1 U7602 ( .A(n1736), .Y(n6472) );
  AND2X1 U7603 ( .A(recentVBools_head_i[30]), .B(n9008), .Y(n1714) );
  INVX1 U7604 ( .A(n1714), .Y(n6473) );
  AND2X1 U7605 ( .A(n2756), .B(n8992), .Y(n1621) );
  INVX1 U7606 ( .A(n1621), .Y(n6474) );
  BUFX2 U7607 ( .A(n2789), .Y(n6475) );
  BUFX2 U7608 ( .A(n2847), .Y(n6476) );
  BUFX2 U7609 ( .A(n2811), .Y(n6477) );
  BUFX2 U7610 ( .A(n2743), .Y(n6478) );
  AND2X1 U7611 ( .A(CircularBuffer_len_write_assig_fu_817_p2[1]), .B(n1646), 
        .Y(n1601) );
  INVX1 U7612 ( .A(n1601), .Y(n6479) );
  AND2X1 U7613 ( .A(CircularBuffer_sum_read_assign_reg_1610[4]), .B(n9007), 
        .Y(n1458) );
  INVX1 U7614 ( .A(n1458), .Y(n6480) );
  AND2X1 U7615 ( .A(CircularBuffer_sum_read_assign_reg_1610[13]), .B(n9006), 
        .Y(n1440) );
  INVX1 U7616 ( .A(n1440), .Y(n6481) );
  AND2X1 U7617 ( .A(n9012), .B(sum_phi_fu_311_p4[7]), .Y(n2668) );
  INVX1 U7618 ( .A(n2668), .Y(n6482) );
  BUFX2 U7619 ( .A(n2723), .Y(n6483) );
  AND2X1 U7620 ( .A(n9012), .B(sum_phi_fu_311_p4[21]), .Y(n2612) );
  INVX1 U7621 ( .A(n2612), .Y(n6484) );
  BUFX2 U7622 ( .A(n2711), .Y(n6485) );
  AND2X1 U7623 ( .A(recentABools_head_i[5]), .B(n9037), .Y(n1331) );
  INVX1 U7624 ( .A(n1331), .Y(n6486) );
  AND2X1 U7625 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[15]), .B(n9040), 
        .Y(n1309) );
  INVX1 U7626 ( .A(n1309), .Y(n6487) );
  AND2X1 U7627 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[20]), .B(n9039), 
        .Y(n1298) );
  INVX1 U7628 ( .A(n1298), .Y(n6488) );
  AND2X1 U7629 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[26]), .B(n9038), 
        .Y(n1282) );
  INVX1 U7630 ( .A(n1282), .Y(n6489) );
  AND2X1 U7631 ( .A(VbeatFallDelay_new_1_reg_342[4]), .B(n9013), .Y(n2161) );
  INVX1 U7632 ( .A(n2161), .Y(n6490) );
  AND2X1 U7633 ( .A(VbeatFallDelay[5]), .B(n9036), .Y(n1186) );
  INVX1 U7634 ( .A(n1186), .Y(n6491) );
  AND2X1 U7635 ( .A(tmp_5_fu_726_p2[9]), .B(n8993), .Y(n1172) );
  INVX1 U7636 ( .A(n1172), .Y(n6492) );
  AND2X1 U7637 ( .A(VbeatFallDelay[16]), .B(n9035), .Y(n1142) );
  INVX1 U7638 ( .A(n1142), .Y(n6493) );
  AND2X1 U7639 ( .A(VbeatFallDelay_new_1_reg_342[18]), .B(n9013), .Y(n2175) );
  INVX1 U7640 ( .A(n2175), .Y(n6494) );
  AND2X1 U7641 ( .A(tmp_5_fu_726_p2[26]), .B(n8994), .Y(n1104) );
  INVX1 U7642 ( .A(n1104), .Y(n6495) );
  AND2X1 U7643 ( .A(VbeatFallDelay[27]), .B(n9034), .Y(n1098) );
  INVX1 U7644 ( .A(n1098), .Y(n6496) );
  AND2X1 U7645 ( .A(VbeatDelay[2]), .B(n9033), .Y(n1069) );
  INVX1 U7646 ( .A(n1069), .Y(n6497) );
  AND2X1 U7647 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[10]), .Y(n2556) );
  INVX1 U7648 ( .A(n2556), .Y(n6498) );
  AND2X1 U7649 ( .A(tmp_4_fu_716_p2[13]), .B(n8995), .Y(n1036) );
  INVX1 U7650 ( .A(n1036), .Y(n6499) );
  AND2X1 U7651 ( .A(VbeatDelay[15]), .B(n9032), .Y(n1028) );
  INVX1 U7652 ( .A(n1028), .Y(n6500) );
  AND2X1 U7653 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[21]), .Y(n2545) );
  INVX1 U7654 ( .A(n2545), .Y(n6501) );
  AND2X1 U7655 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[3]), .Y(n2418) );
  INVX1 U7656 ( .A(n2418), .Y(n6502) );
  BUFX2 U7657 ( .A(n2328), .Y(n6503) );
  AND2X1 U7658 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[10]), .Y(n2446) );
  INVX1 U7659 ( .A(n2446), .Y(n6504) );
  BUFX2 U7660 ( .A(n2311), .Y(n6505) );
  AND2X1 U7661 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[23]), .Y(n2498) );
  INVX1 U7662 ( .A(n2498), .Y(n6506) );
  AND2X1 U7663 ( .A(n2285), .B(n9019), .Y(n961) );
  INVX1 U7664 ( .A(n961), .Y(n6507) );
  BUFX2 U7665 ( .A(n2392), .Y(n6508) );
  BUFX2 U7666 ( .A(n2290), .Y(n6509) );
  BUFX2 U7667 ( .A(n2366), .Y(n6510) );
  AND2X1 U7668 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[1]), .B(n970), 
        .Y(n925) );
  INVX1 U7669 ( .A(n925), .Y(n6511) );
  AND2X1 U7670 ( .A(AbeatDelay_new_reg_394[0]), .B(n9041), .Y(n2234) );
  INVX1 U7671 ( .A(n2234), .Y(n6512) );
  AND2X1 U7672 ( .A(tmp_3_fu_706_p2[1]), .B(n8996), .Y(n790) );
  INVX1 U7673 ( .A(n790), .Y(n6513) );
  AND2X1 U7674 ( .A(AbeatDelay[9]), .B(n8896), .Y(n761) );
  INVX1 U7675 ( .A(n761), .Y(n6514) );
  AND2X1 U7676 ( .A(tmp_3_fu_706_p2[19]), .B(n8997), .Y(n729) );
  INVX1 U7677 ( .A(n729), .Y(n6515) );
  AND2X1 U7678 ( .A(AbeatDelay_new_reg_394[20]), .B(n9041), .Y(n2214) );
  INVX1 U7679 ( .A(n2214), .Y(n6516) );
  AND2X1 U7680 ( .A(AbeatDelay[28]), .B(n10670), .Y(n696) );
  INVX1 U7681 ( .A(n696), .Y(n6517) );
  AND2X1 U7682 ( .A(AstimDelay[12]), .B(n8896), .Y(n647) );
  INVX1 U7683 ( .A(n647), .Y(n6518) );
  AND2X1 U7684 ( .A(tmp_6_fu_497_p3[14]), .B(n8966), .Y(n642) );
  INVX1 U7685 ( .A(n642), .Y(n6519) );
  AND2X1 U7686 ( .A(AstimDelay[29]), .B(n8896), .Y(n596) );
  INVX1 U7687 ( .A(n596), .Y(n6520) );
  AND2X1 U7688 ( .A(tmp_7_fu_511_p3[2]), .B(n8965), .Y(n578) );
  INVX1 U7689 ( .A(n578), .Y(n6521) );
  AND2X1 U7690 ( .A(VstimDelay[15]), .B(n8896), .Y(n538) );
  INVX1 U7691 ( .A(n538), .Y(n6522) );
  AND2X1 U7692 ( .A(tmp_7_fu_511_p3[18]), .B(n8964), .Y(n530) );
  INVX1 U7693 ( .A(n530), .Y(n6523) );
  AND2X1 U7694 ( .A(\Decision_AXILiteS_s_axi_U/n564 ), .B(
        \Decision_AXILiteS_s_axi_U/n351 ), .Y(\Decision_AXILiteS_s_axi_U/n369 ) );
  INVX1 U7695 ( .A(\Decision_AXILiteS_s_axi_U/n369 ), .Y(n6524) );
  AND2X1 U7696 ( .A(\Decision_AXILiteS_s_axi_U/n366 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n414 ) );
  INVX1 U7697 ( .A(\Decision_AXILiteS_s_axi_U/n414 ), .Y(n6525) );
  AND2X1 U7698 ( .A(\Decision_AXILiteS_s_axi_U/n360 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n453 ) );
  INVX1 U7699 ( .A(\Decision_AXILiteS_s_axi_U/n453 ), .Y(n6526) );
  AND2X1 U7700 ( .A(a_length[25]), .B(n8116), .Y(
        \Decision_AXILiteS_s_axi_U/n427 ) );
  INVX1 U7701 ( .A(\Decision_AXILiteS_s_axi_U/n427 ), .Y(n6527) );
  AND2X1 U7702 ( .A(\Decision_AXILiteS_s_axi_U/n362 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n517 ) );
  INVX1 U7703 ( .A(\Decision_AXILiteS_s_axi_U/n517 ), .Y(n6528) );
  AND2X1 U7704 ( .A(vthresh[24]), .B(n7865), .Y(
        \Decision_AXILiteS_s_axi_U/n491 ) );
  INVX1 U7705 ( .A(\Decision_AXILiteS_s_axi_U/n491 ), .Y(n6529) );
  AND2X1 U7706 ( .A(\Decision_AXILiteS_s_axi_U/n364 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n560 ) );
  INVX1 U7707 ( .A(\Decision_AXILiteS_s_axi_U/n560 ), .Y(n6530) );
  AND2X1 U7708 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[13]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n405 )
         );
  INVX1 U7709 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n405 ), 
        .Y(n6531) );
  AND2X1 U7710 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][15] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n581 )
         );
  INVX1 U7711 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n581 ), 
        .Y(n6532) );
  AND2X1 U7712 ( .A(n9468), .B(data_read_reg_1495[6]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n596 )
         );
  INVX1 U7713 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n596 ), 
        .Y(n6533) );
  AND2X1 U7714 ( .A(n9469), .B(data_read_reg_1495[7]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n632 )
         );
  INVX1 U7715 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n632 ), 
        .Y(n6534) );
  AND2X1 U7716 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][0] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n653 )
         );
  INVX1 U7717 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n653 ), 
        .Y(n6535) );
  AND2X1 U7718 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][12] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n665 )
         );
  INVX1 U7719 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n665 ), 
        .Y(n6536) );
  AND2X1 U7720 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][1] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n673 )
         );
  INVX1 U7721 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n673 ), 
        .Y(n6537) );
  AND2X1 U7722 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][13] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n685 )
         );
  INVX1 U7723 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n685 ), 
        .Y(n6538) );
  AND2X1 U7724 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][2] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n692 )
         );
  INVX1 U7725 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n692 ), 
        .Y(n6539) );
  AND2X1 U7726 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][3] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n710 )
         );
  INVX1 U7727 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n710 ), 
        .Y(n6540) );
  AND2X1 U7728 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][6] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n764 )
         );
  INVX1 U7729 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n764 ), 
        .Y(n6541) );
  AND2X1 U7730 ( .A(n9466), .B(data_read_reg_1495[0]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n776 )
         );
  INVX1 U7731 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n776 ), 
        .Y(n6542) );
  AND2X1 U7732 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][7] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n816 )
         );
  INVX1 U7733 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n816 ), 
        .Y(n6543) );
  AND2X1 U7734 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][4] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n831 )
         );
  INVX1 U7735 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n831 ), 
        .Y(n6544) );
  AND2X1 U7736 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][5] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n849 )
         );
  INVX1 U7737 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n849 ), 
        .Y(n6545) );
  AND2X1 U7738 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[1]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n864 )
         );
  INVX1 U7739 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n864 ), 
        .Y(n6546) );
  AND2X1 U7740 ( .A(sum_reg_308[1]), .B(n8929), .Y(n2694) );
  INVX1 U7741 ( .A(n2694), .Y(n6547) );
  AND2X1 U7742 ( .A(sum_1_reg_376[31]), .B(n8930), .Y(n2532) );
  INVX1 U7743 ( .A(n2532), .Y(n6548) );
  AND2X1 U7744 ( .A(sum_reg_308[12]), .B(n8929), .Y(n2650) );
  INVX1 U7745 ( .A(n2650), .Y(n6549) );
  AND2X1 U7746 ( .A(sum_1_reg_376[13]), .B(n8930), .Y(n2460) );
  INVX1 U7747 ( .A(n2460), .Y(n6550) );
  AND2X1 U7748 ( .A(tmp_29_i_fu_752_p2[28]), .B(n8920), .Y(n3164) );
  INVX1 U7749 ( .A(n3164), .Y(n6551) );
  AND2X1 U7750 ( .A(tmp_29_i1_fu_1065_p2[28]), .B(n8922), .Y(n3216) );
  INVX1 U7751 ( .A(n3216), .Y(n6552) );
  AND2X1 U7752 ( .A(tmp_29_i_fu_752_p2[11]), .B(n8920), .Y(n3182) );
  INVX1 U7753 ( .A(n3182), .Y(n6553) );
  AND2X1 U7754 ( .A(tmp_29_i1_fu_1065_p2[11]), .B(n8922), .Y(n3234) );
  INVX1 U7755 ( .A(n3234), .Y(n6554) );
  AND2X1 U7756 ( .A(n8402), .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n27 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n26 ) );
  INVX1 U7757 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n26 ), 
        .Y(n6555) );
  AND2X1 U7758 ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n119 ), .B(
        recentABools_data_address0[2]), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n29 ) );
  INVX1 U7759 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n29 ), 
        .Y(n6556) );
  INVX1 U7760 ( .A(n4627), .Y(n6557) );
  AND2X1 U7761 ( .A(ACaptureThresh_loc_reg_288[7]), .B(n8971), .Y(n3048) );
  INVX1 U7762 ( .A(n3048), .Y(n6558) );
  BUFX2 U7763 ( .A(n3047), .Y(n6559) );
  INVX1 U7764 ( .A(n4611), .Y(n6560) );
  AND2X1 U7765 ( .A(ACaptureThresh_loc_reg_288[23]), .B(n8971), .Y(n3016) );
  INVX1 U7766 ( .A(n3016), .Y(n6561) );
  BUFX2 U7767 ( .A(n3015), .Y(n6562) );
  INVX1 U7768 ( .A(n4565), .Y(n6563) );
  AND2X1 U7769 ( .A(VCaptureThresh_loc_reg_298[5]), .B(n8970), .Y(n2924) );
  INVX1 U7770 ( .A(n2924), .Y(n6564) );
  BUFX2 U7771 ( .A(n2923), .Y(n6565) );
  INVX1 U7772 ( .A(n4549), .Y(n6566) );
  AND2X1 U7773 ( .A(VCaptureThresh_loc_reg_298[21]), .B(n8969), .Y(n2892) );
  INVX1 U7774 ( .A(n2892), .Y(n6567) );
  BUFX2 U7775 ( .A(n2891), .Y(n6568) );
  AND2X1 U7776 ( .A(recentdatapoints_len_load_op_fu_556_p2[1]), .B(n8972), .Y(
        n2024) );
  INVX1 U7777 ( .A(n2024), .Y(n6569) );
  AND2X1 U7778 ( .A(recentdatapoints_len_load_op_fu_556_p2[17]), .B(n8972), 
        .Y(n1839) );
  INVX1 U7779 ( .A(n1839), .Y(n6570) );
  AND2X1 U7780 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[6]), 
        .Y(n448) );
  INVX1 U7781 ( .A(n448), .Y(n6571) );
  AND2X1 U7782 ( .A(CircularBuffer_len_read_assign_fu_772_p2[24]), .B(n8919), 
        .Y(n2746) );
  INVX1 U7783 ( .A(n2746), .Y(n6572) );
  AND2X1 U7784 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[24]), .B(n8921), .Y(n2253) );
  INVX1 U7785 ( .A(n2253), .Y(n6573) );
  AND2X1 U7786 ( .A(a_flip[7]), .B(n8951), .Y(n3139) );
  INVX1 U7787 ( .A(n3139), .Y(n6574) );
  AND2X1 U7788 ( .A(a_length[2]), .B(n8952), .Y(n3122) );
  INVX1 U7789 ( .A(n3122), .Y(n6575) );
  AND2X1 U7790 ( .A(a_length[23]), .B(n8953), .Y(n3080) );
  INVX1 U7791 ( .A(n3080), .Y(n6576) );
  AND2X1 U7792 ( .A(v_length[15]), .B(n8955), .Y(n2968) );
  INVX1 U7793 ( .A(n2968), .Y(n6577) );
  AND2X1 U7794 ( .A(v_length[25]), .B(n8954), .Y(n2948) );
  INVX1 U7795 ( .A(n2948), .Y(n6578) );
  AND2X1 U7796 ( .A(recentdatapoints_head_i[30]), .B(n8979), .Y(n1953) );
  INVX1 U7797 ( .A(n1953), .Y(n6579) );
  AND2X1 U7798 ( .A(p_tmp_i_reg_1556[27]), .B(n8978), .Y(n1916) );
  INVX1 U7799 ( .A(n1916), .Y(n6580) );
  AND2X1 U7800 ( .A(p_tmp_i_reg_1556[15]), .B(n8980), .Y(n1892) );
  INVX1 U7801 ( .A(n1892), .Y(n6581) );
  AND2X1 U7802 ( .A(CircularBuffer_head_i_read_ass_reg_1624[9]), .B(n9011), 
        .Y(n1778) );
  INVX1 U7803 ( .A(n1778), .Y(n6582) );
  AND2X1 U7804 ( .A(recentVBools_head_i[16]), .B(n9010), .Y(n1756) );
  INVX1 U7805 ( .A(n1756), .Y(n6583) );
  AND2X1 U7806 ( .A(recentVBools_head_i[23]), .B(n9009), .Y(n1735) );
  INVX1 U7807 ( .A(n1735), .Y(n6584) );
  AND2X1 U7808 ( .A(n2742), .B(n8991), .Y(n1610) );
  INVX1 U7809 ( .A(n1610), .Y(n6585) );
  BUFX2 U7810 ( .A(n2845), .Y(n6586) );
  BUFX2 U7811 ( .A(n2775), .Y(n6587) );
  BUFX2 U7812 ( .A(n2749), .Y(n6588) );
  BUFX2 U7813 ( .A(n2809), .Y(n6589) );
  AND2X1 U7814 ( .A(CircularBuffer_len_write_assig_fu_817_p2[2]), .B(n1646), 
        .Y(n1600) );
  INVX1 U7815 ( .A(n1600), .Y(n6590) );
  AND2X1 U7816 ( .A(CircularBuffer_sum_read_assign_reg_1610[5]), .B(n9007), 
        .Y(n1456) );
  INVX1 U7817 ( .A(n1456), .Y(n6591) );
  AND2X1 U7818 ( .A(CircularBuffer_sum_read_assign_reg_1610[14]), .B(n9006), 
        .Y(n1438) );
  INVX1 U7819 ( .A(n1438), .Y(n6592) );
  BUFX2 U7820 ( .A(n2724), .Y(n6593) );
  AND2X1 U7821 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[9]), .Y(n2660) );
  INVX1 U7822 ( .A(n2660), .Y(n6594) );
  AND2X1 U7823 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[22]), .Y(n2608) );
  INVX1 U7824 ( .A(n2608), .Y(n6595) );
  BUFX2 U7825 ( .A(n2710), .Y(n6596) );
  AND2X1 U7826 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[12]), .B(n9034), 
        .Y(n1364) );
  INVX1 U7827 ( .A(n1364), .Y(n6597) );
  AND2X1 U7828 ( .A(recentABools_head_i[18]), .B(n9039), .Y(n1302) );
  INVX1 U7829 ( .A(n1302), .Y(n6598) );
  AND2X1 U7830 ( .A(recentABools_head_i[24]), .B(n9038), .Y(n1286) );
  INVX1 U7831 ( .A(n1286), .Y(n6599) );
  AND2X1 U7832 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[30]), .B(n9037), 
        .Y(n1273) );
  INVX1 U7833 ( .A(n1273), .Y(n6600) );
  AND2X1 U7834 ( .A(tmp_5_fu_726_p2[2]), .B(n8992), .Y(n1200) );
  INVX1 U7835 ( .A(n1200), .Y(n6601) );
  AND2X1 U7836 ( .A(VbeatFallDelay_new_1_reg_342[5]), .B(n9013), .Y(n2162) );
  INVX1 U7837 ( .A(n2162), .Y(n6602) );
  AND2X1 U7838 ( .A(VbeatFallDelay[6]), .B(n9036), .Y(n1182) );
  INVX1 U7839 ( .A(n1182), .Y(n6603) );
  AND2X1 U7840 ( .A(tmp_5_fu_726_p2[10]), .B(n8993), .Y(n1168) );
  INVX1 U7841 ( .A(n1168), .Y(n6604) );
  AND2X1 U7842 ( .A(VbeatFallDelay[17]), .B(n9035), .Y(n1138) );
  INVX1 U7843 ( .A(n1138), .Y(n6605) );
  AND2X1 U7844 ( .A(VbeatFallDelay_new_1_reg_342[19]), .B(n9013), .Y(n2176) );
  INVX1 U7845 ( .A(n2176), .Y(n6606) );
  AND2X1 U7846 ( .A(tmp_5_fu_726_p2[27]), .B(n8994), .Y(n1100) );
  INVX1 U7847 ( .A(n1100), .Y(n6607) );
  AND2X1 U7848 ( .A(VbeatDelay[3]), .B(n9033), .Y(n1080) );
  INVX1 U7849 ( .A(n1080), .Y(n6608) );
  AND2X1 U7850 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[9]), .Y(n2557) );
  INVX1 U7851 ( .A(n2557), .Y(n6609) );
  AND2X1 U7852 ( .A(VbeatDelay[10]), .B(n9032), .Y(n1045) );
  INVX1 U7853 ( .A(n1045), .Y(n6610) );
  AND2X1 U7854 ( .A(tmp_4_fu_716_p2[14]), .B(n8995), .Y(n1033) );
  INVX1 U7855 ( .A(n1033), .Y(n6611) );
  AND2X1 U7856 ( .A(VbeatDelay[16]), .B(n9031), .Y(n1025) );
  INVX1 U7857 ( .A(n1025), .Y(n6612) );
  AND2X1 U7858 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[22]), .Y(n2544) );
  INVX1 U7859 ( .A(n2544), .Y(n6613) );
  BUFX2 U7860 ( .A(n2334), .Y(n6614) );
  AND2X1 U7861 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[2]), .Y(n2414) );
  INVX1 U7862 ( .A(n2414), .Y(n6615) );
  AND2X1 U7863 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[12]), .Y(n2454) );
  INVX1 U7864 ( .A(n2454), .Y(n6616) );
  BUFX2 U7865 ( .A(n2321), .Y(n6617) );
  AND2X1 U7866 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[24]), .Y(n2502) );
  INVX1 U7867 ( .A(n2502), .Y(n6618) );
  BUFX2 U7868 ( .A(n2307), .Y(n6619) );
  BUFX2 U7869 ( .A(n2390), .Y(n6620) );
  BUFX2 U7870 ( .A(n2288), .Y(n6621) );
  BUFX2 U7871 ( .A(n2364), .Y(n6622) );
  AND2X1 U7872 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[2]), .B(n970), 
        .Y(n924) );
  INVX1 U7873 ( .A(n924), .Y(n6623) );
  AND2X1 U7874 ( .A(n10671), .B(n8996), .Y(n792) );
  INVX1 U7875 ( .A(n792), .Y(n6624) );
  AND2X1 U7876 ( .A(AbeatDelay_new_reg_394[1]), .B(n9041), .Y(n2233) );
  INVX1 U7877 ( .A(n2233), .Y(n6625) );
  AND2X1 U7878 ( .A(AbeatDelay[15]), .B(n8896), .Y(n741) );
  INVX1 U7879 ( .A(n741), .Y(n6626) );
  AND2X1 U7880 ( .A(tmp_3_fu_706_p2[20]), .B(n8997), .Y(n725) );
  INVX1 U7881 ( .A(n725), .Y(n6627) );
  AND2X1 U7882 ( .A(AbeatDelay_new_reg_394[21]), .B(n9041), .Y(n2213) );
  INVX1 U7883 ( .A(n2213), .Y(n6628) );
  AND2X1 U7884 ( .A(AbeatDelay[29]), .B(n8896), .Y(n692) );
  INVX1 U7885 ( .A(n692), .Y(n6629) );
  AND2X1 U7886 ( .A(n10742), .B(n8967), .Y(n683) );
  INVX1 U7887 ( .A(n683), .Y(n6630) );
  AND2X1 U7888 ( .A(AstimDelay[13]), .B(n8896), .Y(n644) );
  INVX1 U7889 ( .A(n644), .Y(n6631) );
  AND2X1 U7890 ( .A(tmp_6_fu_497_p3[15]), .B(n8966), .Y(n639) );
  INVX1 U7891 ( .A(n639), .Y(n6632) );
  AND2X1 U7892 ( .A(AstimDelay[30]), .B(n10670), .Y(n593) );
  INVX1 U7893 ( .A(n593), .Y(n6633) );
  AND2X1 U7894 ( .A(tmp_7_fu_511_p3[3]), .B(n8965), .Y(n575) );
  INVX1 U7895 ( .A(n575), .Y(n6634) );
  AND2X1 U7896 ( .A(VstimDelay[16]), .B(n8896), .Y(n535) );
  INVX1 U7897 ( .A(n535), .Y(n6635) );
  AND2X1 U7898 ( .A(tmp_7_fu_511_p3[19]), .B(n8964), .Y(n527) );
  INVX1 U7899 ( .A(n527), .Y(n6636) );
  AND2X1 U7900 ( .A(\Decision_AXILiteS_s_axi_U/n368 ), .B(
        \Decision_AXILiteS_s_axi_U/n351 ), .Y(\Decision_AXILiteS_s_axi_U/n367 ) );
  INVX1 U7901 ( .A(\Decision_AXILiteS_s_axi_U/n367 ), .Y(n6637) );
  AND2X1 U7902 ( .A(\Decision_AXILiteS_s_axi_U/n358 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n410 ) );
  INVX1 U7903 ( .A(\Decision_AXILiteS_s_axi_U/n410 ), .Y(n6638) );
  AND2X1 U7904 ( .A(\Decision_AXILiteS_s_axi_U/n364 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n455 ) );
  INVX1 U7905 ( .A(\Decision_AXILiteS_s_axi_U/n455 ), .Y(n6639) );
  AND2X1 U7906 ( .A(\Decision_AXILiteS_s_axi_U/n360 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n516 ) );
  INVX1 U7907 ( .A(\Decision_AXILiteS_s_axi_U/n516 ), .Y(n6640) );
  AND2X1 U7908 ( .A(vthresh[25]), .B(n7865), .Y(
        \Decision_AXILiteS_s_axi_U/n490 ) );
  INVX1 U7909 ( .A(\Decision_AXILiteS_s_axi_U/n490 ), .Y(n6641) );
  AND2X1 U7910 ( .A(\Decision_AXILiteS_s_axi_U/n362 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n559 ) );
  INVX1 U7911 ( .A(\Decision_AXILiteS_s_axi_U/n559 ), .Y(n6642) );
  AND2X1 U7912 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[14]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n407 )
         );
  INVX1 U7913 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n407 ), 
        .Y(n6643) );
  AND2X1 U7914 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][0] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n551 )
         );
  INVX1 U7915 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n551 ), 
        .Y(n6644) );
  AND2X1 U7916 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][12] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n575 )
         );
  INVX1 U7917 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n575 ), 
        .Y(n6645) );
  AND2X1 U7918 ( .A(n9468), .B(data_read_reg_1495[1]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n586 )
         );
  INVX1 U7919 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n586 ), 
        .Y(n6646) );
  AND2X1 U7920 ( .A(n9469), .B(data_read_reg_1495[0]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n618 )
         );
  INVX1 U7921 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n618 ), 
        .Y(n6647) );
  AND2X1 U7922 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][15] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n668 )
         );
  INVX1 U7923 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n668 ), 
        .Y(n6648) );
  AND2X1 U7924 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][14] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n686 )
         );
  INVX1 U7925 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n686 ), 
        .Y(n6649) );
  AND2X1 U7926 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][3] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n727 )
         );
  INVX1 U7927 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n727 ), 
        .Y(n6650) );
  AND2X1 U7928 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][2] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n743 )
         );
  INVX1 U7929 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n743 ), 
        .Y(n6651) );
  AND2X1 U7930 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][5] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n763 )
         );
  INVX1 U7931 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n763 ), 
        .Y(n6652) );
  AND2X1 U7932 ( .A(n9466), .B(data_read_reg_1495[7]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n790 )
         );
  INVX1 U7933 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n790 ), 
        .Y(n6653) );
  AND2X1 U7934 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][4] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n813 )
         );
  INVX1 U7935 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n813 ), 
        .Y(n6654) );
  AND2X1 U7936 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][7] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n834 )
         );
  INVX1 U7937 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n834 ), 
        .Y(n6655) );
  AND2X1 U7938 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][6] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n850 )
         );
  INVX1 U7939 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n850 ), 
        .Y(n6656) );
  AND2X1 U7940 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[6]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n874 )
         );
  INVX1 U7941 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n874 ), 
        .Y(n6657) );
  AND2X1 U7942 ( .A(sum_reg_308[28]), .B(n8929), .Y(n2586) );
  INVX1 U7943 ( .A(n2586), .Y(n6658) );
  AND2X1 U7944 ( .A(sum_1_reg_376[3]), .B(n8930), .Y(n2420) );
  INVX1 U7945 ( .A(n2420), .Y(n6659) );
  AND2X1 U7946 ( .A(sum_reg_308[4]), .B(n8929), .Y(n2682) );
  INVX1 U7947 ( .A(n2682), .Y(n6660) );
  AND2X1 U7948 ( .A(sum_1_reg_376[16]), .B(n8930), .Y(n2472) );
  INVX1 U7949 ( .A(n2472), .Y(n6661) );
  AND2X1 U7950 ( .A(tmp_29_i_fu_752_p2[20]), .B(n8920), .Y(n3172) );
  INVX1 U7951 ( .A(n3172), .Y(n6662) );
  AND2X1 U7952 ( .A(tmp_29_i1_fu_1065_p2[20]), .B(n8922), .Y(n3224) );
  INVX1 U7953 ( .A(n3224), .Y(n6663) );
  AND2X1 U7954 ( .A(tmp_29_i_fu_752_p2[10]), .B(n8920), .Y(n3183) );
  INVX1 U7955 ( .A(n3183), .Y(n6664) );
  AND2X1 U7956 ( .A(tmp_29_i1_fu_1065_p2[10]), .B(n8922), .Y(n3235) );
  INVX1 U7957 ( .A(n3235), .Y(n6665) );
  INVX1 U7958 ( .A(n4626), .Y(n6666) );
  AND2X1 U7959 ( .A(ACaptureThresh_loc_reg_288[8]), .B(n8968), .Y(n3046) );
  INVX1 U7960 ( .A(n3046), .Y(n6667) );
  BUFX2 U7961 ( .A(n3045), .Y(n6668) );
  INVX1 U7962 ( .A(n4610), .Y(n6669) );
  AND2X1 U7963 ( .A(ACaptureThresh_loc_reg_288[24]), .B(n8971), .Y(n3014) );
  INVX1 U7964 ( .A(n3014), .Y(n6670) );
  BUFX2 U7965 ( .A(n3013), .Y(n6671) );
  INVX1 U7966 ( .A(n4563), .Y(n6672) );
  AND2X1 U7967 ( .A(VCaptureThresh_loc_reg_298[7]), .B(n8970), .Y(n2920) );
  INVX1 U7968 ( .A(n2920), .Y(n6673) );
  BUFX2 U7969 ( .A(n2919), .Y(n6674) );
  INVX1 U7970 ( .A(n4548), .Y(n6675) );
  AND2X1 U7971 ( .A(VCaptureThresh_loc_reg_298[22]), .B(n8969), .Y(n2890) );
  INVX1 U7972 ( .A(n2890), .Y(n6676) );
  BUFX2 U7973 ( .A(n2889), .Y(n6677) );
  BUFX2 U7974 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n31 ), 
        .Y(n6678) );
  BUFX2 U7975 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n32 ), 
        .Y(n6679) );
  BUFX2 U7976 ( .A(n1801), .Y(n6680) );
  BUFX2 U7977 ( .A(n1802), .Y(n6681) );
  BUFX2 U7978 ( .A(n1231), .Y(n6682) );
  BUFX2 U7979 ( .A(n1232), .Y(n6683) );
  AND2X1 U7980 ( .A(recentdatapoints_len_load_op_fu_556_p2[3]), .B(n8972), .Y(
        n1823) );
  INVX1 U7981 ( .A(n1823), .Y(n6684) );
  AND2X1 U7982 ( .A(recentdatapoints_len_load_op_fu_556_p2[18]), .B(n8972), 
        .Y(n1840) );
  INVX1 U7983 ( .A(n1840), .Y(n6685) );
  AND2X1 U7984 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[11]), 
        .Y(n467) );
  INVX1 U7985 ( .A(n467), .Y(n6686) );
  AND2X1 U7986 ( .A(CircularBuffer_len_read_assign_fu_772_p2[28]), .B(n8919), 
        .Y(n2738) );
  INVX1 U7987 ( .A(n2738), .Y(n6687) );
  AND2X1 U7988 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[28]), .B(n8921), .Y(n2245) );
  INVX1 U7989 ( .A(n2245), .Y(n6688) );
  AND2X1 U7990 ( .A(v_flip[1]), .B(n8951), .Y(n3136) );
  INVX1 U7991 ( .A(n3136), .Y(n6689) );
  AND2X1 U7992 ( .A(a_length[3]), .B(n8952), .Y(n3120) );
  INVX1 U7993 ( .A(n3120), .Y(n6690) );
  AND2X1 U7994 ( .A(a_length[24]), .B(n8953), .Y(n3078) );
  INVX1 U7995 ( .A(n3078), .Y(n6691) );
  AND2X1 U7996 ( .A(v_length[16]), .B(n8955), .Y(n2966) );
  INVX1 U7997 ( .A(n2966), .Y(n6692) );
  AND2X1 U7998 ( .A(v_length[26]), .B(n8954), .Y(n2946) );
  INVX1 U7999 ( .A(n2946), .Y(n6693) );
  AND2X1 U8000 ( .A(n8963), .B(recentdatapoints_head_i[0]), .Y(n1986) );
  INVX1 U8001 ( .A(n1986), .Y(n6694) );
  AND2X1 U8002 ( .A(p_tmp_i_reg_1556[31]), .B(n8979), .Y(n1924) );
  INVX1 U8003 ( .A(n1924), .Y(n6695) );
  AND2X1 U8004 ( .A(p_tmp_i_reg_1556[21]), .B(n8980), .Y(n1904) );
  INVX1 U8005 ( .A(n1904), .Y(n6696) );
  AND2X1 U8006 ( .A(p_tmp_i_reg_1556[14]), .B(n8980), .Y(n1890) );
  INVX1 U8007 ( .A(n1890), .Y(n6697) );
  AND2X1 U8008 ( .A(recentVBools_head_i[9]), .B(n9011), .Y(n1777) );
  INVX1 U8009 ( .A(n1777), .Y(n6698) );
  AND2X1 U8010 ( .A(CircularBuffer_head_i_read_ass_reg_1624[17]), .B(n9010), 
        .Y(n1754) );
  INVX1 U8011 ( .A(n1754), .Y(n6699) );
  AND2X1 U8012 ( .A(n2740), .B(n8991), .Y(n1609) );
  INVX1 U8013 ( .A(n1609), .Y(n6700) );
  BUFX2 U8014 ( .A(n2787), .Y(n6701) );
  BUFX2 U8015 ( .A(n2843), .Y(n6702) );
  BUFX2 U8016 ( .A(n2773), .Y(n6703) );
  BUFX2 U8017 ( .A(n2745), .Y(n6704) );
  BUFX2 U8018 ( .A(n2807), .Y(n6705) );
  AND2X1 U8019 ( .A(CircularBuffer_len_write_assig_fu_817_p2[3]), .B(n1646), 
        .Y(n1598) );
  INVX1 U8020 ( .A(n1598), .Y(n6706) );
  AND2X1 U8021 ( .A(CircularBuffer_len_write_assig_fu_817_p2[7]), .B(n8894), 
        .Y(n1592) );
  INVX1 U8022 ( .A(n1592), .Y(n6707) );
  AND2X1 U8023 ( .A(CircularBuffer_sum_read_assign_reg_1610[6]), .B(n9007), 
        .Y(n1454) );
  INVX1 U8024 ( .A(n1454), .Y(n6708) );
  AND2X1 U8025 ( .A(CircularBuffer_sum_read_assign_reg_1610[15]), .B(n9006), 
        .Y(n1436) );
  INVX1 U8026 ( .A(n1436), .Y(n6709) );
  AND2X1 U8027 ( .A(n9012), .B(sum_phi_fu_311_p4[8]), .Y(n2664) );
  INVX1 U8028 ( .A(n2664), .Y(n6710) );
  BUFX2 U8029 ( .A(n2722), .Y(n6711) );
  AND2X1 U8030 ( .A(n9012), .B(sum_phi_fu_311_p4[23]), .Y(n2604) );
  INVX1 U8031 ( .A(n2604), .Y(n6712) );
  BUFX2 U8032 ( .A(n2708), .Y(n6713) );
  AND2X1 U8033 ( .A(recentABools_head_i[8]), .B(n9038), .Y(n1325) );
  INVX1 U8034 ( .A(n1325), .Y(n6714) );
  AND2X1 U8035 ( .A(recentABools_head_i[15]), .B(n9040), .Y(n1308) );
  INVX1 U8036 ( .A(n1308), .Y(n6715) );
  AND2X1 U8037 ( .A(recentABools_head_i[20]), .B(n9039), .Y(n1297) );
  INVX1 U8038 ( .A(n1297), .Y(n6716) );
  AND2X1 U8039 ( .A(recentABools_head_i[30]), .B(n9037), .Y(n1272) );
  INVX1 U8040 ( .A(n1272), .Y(n6717) );
  AND2X1 U8041 ( .A(tmp_5_fu_726_p2[3]), .B(n8992), .Y(n1196) );
  INVX1 U8042 ( .A(n1196), .Y(n6718) );
  AND2X1 U8043 ( .A(VbeatFallDelay_new_1_reg_342[6]), .B(n9013), .Y(n2163) );
  INVX1 U8044 ( .A(n2163), .Y(n6719) );
  AND2X1 U8045 ( .A(VbeatFallDelay[7]), .B(n9036), .Y(n1178) );
  INVX1 U8046 ( .A(n1178), .Y(n6720) );
  AND2X1 U8047 ( .A(tmp_5_fu_726_p2[8]), .B(n8993), .Y(n1176) );
  INVX1 U8048 ( .A(n1176), .Y(n6721) );
  AND2X1 U8049 ( .A(VbeatFallDelay[18]), .B(n9035), .Y(n1134) );
  INVX1 U8050 ( .A(n1134), .Y(n6722) );
  AND2X1 U8051 ( .A(VbeatFallDelay_new_1_reg_342[20]), .B(n9013), .Y(n2177) );
  INVX1 U8052 ( .A(n2177), .Y(n6723) );
  AND2X1 U8053 ( .A(tmp_5_fu_726_p2[28]), .B(n8994), .Y(n1096) );
  INVX1 U8054 ( .A(n1096), .Y(n6724) );
  AND2X1 U8055 ( .A(VbeatFallDelay[28]), .B(n9034), .Y(n1094) );
  INVX1 U8056 ( .A(n1094), .Y(n6725) );
  AND2X1 U8057 ( .A(VbeatDelay[5]), .B(n9033), .Y(n1060) );
  INVX1 U8058 ( .A(n1060), .Y(n6726) );
  AND2X1 U8059 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[11]), .Y(n2555) );
  INVX1 U8060 ( .A(n2555), .Y(n6727) );
  AND2X1 U8061 ( .A(tmp_4_fu_716_p2[15]), .B(n8995), .Y(n1030) );
  INVX1 U8062 ( .A(n1030), .Y(n6728) );
  AND2X1 U8063 ( .A(VbeatDelay[17]), .B(n9032), .Y(n1021) );
  INVX1 U8064 ( .A(n1021), .Y(n6729) );
  AND2X1 U8065 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[23]), .Y(n2543) );
  INVX1 U8066 ( .A(n2543), .Y(n6730) );
  BUFX2 U8067 ( .A(n2333), .Y(n6731) );
  AND2X1 U8068 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[4]), .Y(n2422) );
  INVX1 U8069 ( .A(n2422), .Y(n6732) );
  AND2X1 U8070 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[13]), .Y(n2458) );
  INVX1 U8071 ( .A(n2458), .Y(n6733) );
  BUFX2 U8072 ( .A(n2320), .Y(n6734) );
  AND2X1 U8073 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[25]), .Y(n2506) );
  INVX1 U8074 ( .A(n2506), .Y(n6735) );
  BUFX2 U8075 ( .A(n2308), .Y(n6736) );
  AND2X1 U8076 ( .A(n2283), .B(n9019), .Y(n959) );
  INVX1 U8077 ( .A(n959), .Y(n6737) );
  BUFX2 U8078 ( .A(n2388), .Y(n6738) );
  BUFX2 U8079 ( .A(n2286), .Y(n6739) );
  BUFX2 U8080 ( .A(n2362), .Y(n6740) );
  AND2X1 U8081 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[3]), .B(n970), 
        .Y(n922) );
  INVX1 U8082 ( .A(n922), .Y(n6741) );
  AND2X1 U8083 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[7]), .B(n8891), 
        .Y(n916) );
  INVX1 U8084 ( .A(n916), .Y(n6742) );
  AND2X1 U8085 ( .A(AbeatDelay[1]), .B(n8896), .Y(n788) );
  INVX1 U8086 ( .A(n788), .Y(n6743) );
  AND2X1 U8087 ( .A(tmp_3_fu_706_p2[3]), .B(n8996), .Y(n783) );
  INVX1 U8088 ( .A(n783), .Y(n6744) );
  AND2X1 U8089 ( .A(AbeatDelay_new_reg_394[7]), .B(n9041), .Y(n2227) );
  INVX1 U8090 ( .A(n2227), .Y(n6745) );
  AND2X1 U8091 ( .A(AbeatDelay[16]), .B(n10670), .Y(n737) );
  INVX1 U8092 ( .A(n737), .Y(n6746) );
  AND2X1 U8093 ( .A(tmp_3_fu_706_p2[21]), .B(n8997), .Y(n722) );
  INVX1 U8094 ( .A(n722), .Y(n6747) );
  AND2X1 U8095 ( .A(AbeatDelay_new_reg_394[22]), .B(n9041), .Y(n2212) );
  INVX1 U8096 ( .A(n2212), .Y(n6748) );
  AND2X1 U8097 ( .A(tmp_6_fu_497_p3[1]), .B(n8967), .Y(n681) );
  INVX1 U8098 ( .A(n681), .Y(n6749) );
  AND2X1 U8099 ( .A(AstimDelay[14]), .B(n8896), .Y(n641) );
  INVX1 U8100 ( .A(n641), .Y(n6750) );
  AND2X1 U8101 ( .A(tmp_6_fu_497_p3[16]), .B(n8966), .Y(n636) );
  INVX1 U8102 ( .A(n636), .Y(n6751) );
  AND2X1 U8103 ( .A(AstimDelay[31]), .B(n8896), .Y(n588) );
  INVX1 U8104 ( .A(n588), .Y(n6752) );
  AND2X1 U8105 ( .A(VstimDelay[0]), .B(n10670), .Y(n584) );
  INVX1 U8106 ( .A(n584), .Y(n6753) );
  AND2X1 U8107 ( .A(tmp_7_fu_511_p3[4]), .B(n8965), .Y(n572) );
  INVX1 U8108 ( .A(n572), .Y(n6754) );
  AND2X1 U8109 ( .A(VstimDelay[17]), .B(n10670), .Y(n532) );
  INVX1 U8110 ( .A(n532), .Y(n6755) );
  AND2X1 U8111 ( .A(tmp_7_fu_511_p3[20]), .B(n8964), .Y(n524) );
  INVX1 U8112 ( .A(n524), .Y(n6756) );
  AND2X1 U8113 ( .A(\Decision_AXILiteS_s_axi_U/n366 ), .B(
        \Decision_AXILiteS_s_axi_U/n351 ), .Y(\Decision_AXILiteS_s_axi_U/n365 ) );
  INVX1 U8114 ( .A(\Decision_AXILiteS_s_axi_U/n365 ), .Y(n6757) );
  AND2X1 U8115 ( .A(\Decision_AXILiteS_s_axi_U/n362 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n454 ) );
  INVX1 U8116 ( .A(\Decision_AXILiteS_s_axi_U/n454 ), .Y(n6758) );
  AND2X1 U8117 ( .A(a_length[27]), .B(n8116), .Y(
        \Decision_AXILiteS_s_axi_U/n425 ) );
  INVX1 U8118 ( .A(\Decision_AXILiteS_s_axi_U/n425 ), .Y(n6759) );
  AND2X1 U8119 ( .A(\Decision_AXILiteS_s_axi_U/n564 ), .B(n8411), .Y(
        \Decision_AXILiteS_s_axi_U/n469 ) );
  INVX1 U8120 ( .A(\Decision_AXILiteS_s_axi_U/n469 ), .Y(n6760) );
  AND2X1 U8121 ( .A(vthresh[26]), .B(n7865), .Y(
        \Decision_AXILiteS_s_axi_U/n489 ) );
  INVX1 U8122 ( .A(\Decision_AXILiteS_s_axi_U/n489 ), .Y(n6761) );
  AND2X1 U8123 ( .A(\Decision_AXILiteS_s_axi_U/n360 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n558 ) );
  INVX1 U8124 ( .A(\Decision_AXILiteS_s_axi_U/n558 ), .Y(n6762) );
  AND2X1 U8125 ( .A(n8393), .B(\Decision_AXILiteS_s_axi_U/n579 ), .Y(
        \Decision_AXILiteS_s_axi_U/n586 ) );
  INVX1 U8126 ( .A(\Decision_AXILiteS_s_axi_U/n586 ), .Y(n6763) );
  AND2X1 U8127 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[15]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n409 )
         );
  INVX1 U8128 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n409 ), 
        .Y(n6764) );
  AND2X1 U8129 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][1] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n553 )
         );
  INVX1 U8130 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n553 ), 
        .Y(n6765) );
  AND2X1 U8131 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][13] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n577 )
         );
  INVX1 U8132 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n577 ), 
        .Y(n6766) );
  AND2X1 U8133 ( .A(n9468), .B(data_read_reg_1495[0]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n584 )
         );
  INVX1 U8134 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n584 ), 
        .Y(n6767) );
  AND2X1 U8135 ( .A(n9469), .B(data_read_reg_1495[1]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n620 )
         );
  INVX1 U8136 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n620 ), 
        .Y(n6768) );
  AND2X1 U8137 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][14] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n667 )
         );
  INVX1 U8138 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n667 ), 
        .Y(n6769) );
  AND2X1 U8139 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][15] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n687 )
         );
  INVX1 U8140 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n687 ), 
        .Y(n6770) );
  AND2X1 U8141 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][2] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n726 )
         );
  INVX1 U8142 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n726 ), 
        .Y(n6771) );
  AND2X1 U8143 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][3] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n744 )
         );
  INVX1 U8144 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n744 ), 
        .Y(n6772) );
  AND2X1 U8145 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][4] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n762 )
         );
  INVX1 U8146 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n762 ), 
        .Y(n6773) );
  AND2X1 U8147 ( .A(n9466), .B(data_read_reg_1495[6]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n788 )
         );
  INVX1 U8148 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n788 ), 
        .Y(n6774) );
  AND2X1 U8149 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][5] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n814 )
         );
  INVX1 U8150 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n814 ), 
        .Y(n6775) );
  AND2X1 U8151 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][6] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n833 )
         );
  INVX1 U8152 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n833 ), 
        .Y(n6776) );
  AND2X1 U8153 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][7] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n851 )
         );
  INVX1 U8154 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n851 ), 
        .Y(n6777) );
  AND2X1 U8155 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[7]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n876 )
         );
  INVX1 U8156 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n876 ), 
        .Y(n6778) );
  AND2X1 U8157 ( .A(sum_reg_308[13]), .B(n8929), .Y(n2646) );
  INVX1 U8158 ( .A(n2646), .Y(n6779) );
  AND2X1 U8159 ( .A(tmp_29_i_fu_752_p2[27]), .B(n8920), .Y(n3165) );
  INVX1 U8160 ( .A(n3165), .Y(n6780) );
  AND2X1 U8161 ( .A(sum_1_reg_376[20]), .B(n8930), .Y(n2488) );
  INVX1 U8162 ( .A(n2488), .Y(n6781) );
  AND2X1 U8163 ( .A(tmp_29_i1_fu_1065_p2[27]), .B(n8922), .Y(n3217) );
  INVX1 U8164 ( .A(n3217), .Y(n6782) );
  AND2X1 U8165 ( .A(sum_1_reg_376[10]), .B(n8930), .Y(n2448) );
  INVX1 U8166 ( .A(n2448), .Y(n6783) );
  AND2X1 U8167 ( .A(tmp_29_i_fu_752_p2[9]), .B(n8920), .Y(n3153) );
  INVX1 U8168 ( .A(n3153), .Y(n6784) );
  AND2X1 U8169 ( .A(tmp_29_i1_fu_1065_p2[9]), .B(n8922), .Y(n3205) );
  INVX1 U8170 ( .A(n3205), .Y(n6785) );
  AND2X1 U8171 ( .A(sum_reg_308[26]), .B(n8929), .Y(n2594) );
  INVX1 U8172 ( .A(n2594), .Y(n6786) );
  INVX1 U8173 ( .A(n4624), .Y(n6787) );
  AND2X1 U8174 ( .A(ACaptureThresh_loc_reg_288[10]), .B(n8971), .Y(n3042) );
  INVX1 U8175 ( .A(n3042), .Y(n6788) );
  BUFX2 U8176 ( .A(n3041), .Y(n6789) );
  INVX1 U8177 ( .A(n4608), .Y(n6790) );
  AND2X1 U8178 ( .A(ACaptureThresh_loc_reg_288[26]), .B(n8971), .Y(n3010) );
  INVX1 U8179 ( .A(n3010), .Y(n6791) );
  BUFX2 U8180 ( .A(n3009), .Y(n6792) );
  INVX1 U8181 ( .A(n4562), .Y(n6793) );
  AND2X1 U8182 ( .A(VCaptureThresh_loc_reg_298[8]), .B(n8970), .Y(n2918) );
  INVX1 U8183 ( .A(n2918), .Y(n6794) );
  BUFX2 U8184 ( .A(n2917), .Y(n6795) );
  INVX1 U8185 ( .A(n4547), .Y(n6796) );
  AND2X1 U8186 ( .A(VCaptureThresh_loc_reg_298[23]), .B(n8969), .Y(n2888) );
  INVX1 U8187 ( .A(n2888), .Y(n6797) );
  BUFX2 U8188 ( .A(n2887), .Y(n6798) );
  BUFX2 U8189 ( .A(n2052), .Y(n6799) );
  BUFX2 U8190 ( .A(n2051), .Y(n6800) );
  BUFX2 U8191 ( .A(n379), .Y(n6801) );
  BUFX2 U8192 ( .A(n378), .Y(n6802) );
  BUFX2 U8193 ( .A(n393), .Y(n6803) );
  BUFX2 U8194 ( .A(n392), .Y(n6804) );
  AND2X1 U8195 ( .A(n9943), .B(n9942), .Y(n1821) );
  INVX1 U8196 ( .A(n1821), .Y(n6805) );
  AND2X1 U8197 ( .A(n10251), .B(n10250), .Y(n1267) );
  INVX1 U8198 ( .A(n1267), .Y(n6806) );
  AND2X1 U8199 ( .A(n9855), .B(n9856), .Y(n2046) );
  INVX1 U8200 ( .A(n2046), .Y(n6807) );
  AND2X1 U8201 ( .A(recentdatapoints_len_load_op_fu_556_p2[5]), .B(n8972), .Y(
        n1825) );
  INVX1 U8202 ( .A(n1825), .Y(n6808) );
  AND2X1 U8203 ( .A(recentdatapoints_len_load_op_fu_556_p2[19]), .B(n8972), 
        .Y(n1841) );
  INVX1 U8204 ( .A(n1841), .Y(n6809) );
  AND2X1 U8205 ( .A(\Decision_AXILiteS_s_axi_U/waddr[4] ), .B(
        \Decision_AXILiteS_s_axi_U/waddr[3] ), .Y(
        \Decision_AXILiteS_s_axi_U/n417 ) );
  INVX1 U8206 ( .A(\Decision_AXILiteS_s_axi_U/n417 ), .Y(n6810) );
  AND2X1 U8207 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[8]), 
        .Y(n444) );
  INVX1 U8208 ( .A(n444), .Y(n6811) );
  AND2X1 U8209 ( .A(CircularBuffer_len_read_assign_fu_772_p2[26]), .B(n8919), 
        .Y(n2742) );
  INVX1 U8210 ( .A(n2742), .Y(n6812) );
  AND2X1 U8211 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[26]), .B(n8921), .Y(n2249) );
  INVX1 U8212 ( .A(n2249), .Y(n6813) );
  AND2X1 U8213 ( .A(v_flip[5]), .B(n8951), .Y(n3130) );
  INVX1 U8214 ( .A(n3130), .Y(n6814) );
  AND2X1 U8215 ( .A(a_length[9]), .B(n8952), .Y(n3108) );
  INVX1 U8216 ( .A(n3108), .Y(n6815) );
  AND2X1 U8217 ( .A(a_length[25]), .B(n8953), .Y(n3076) );
  INVX1 U8218 ( .A(n3076), .Y(n6816) );
  AND2X1 U8219 ( .A(v_length[17]), .B(n8955), .Y(n2964) );
  INVX1 U8220 ( .A(n2964), .Y(n6817) );
  AND2X1 U8221 ( .A(v_length[27]), .B(n8954), .Y(n2944) );
  INVX1 U8222 ( .A(n2944), .Y(n6818) );
  AND2X1 U8223 ( .A(n8963), .B(recentdatapoints_head_i[1]), .Y(n1983) );
  INVX1 U8224 ( .A(n1983), .Y(n6819) );
  AND2X1 U8225 ( .A(recentdatapoints_head_i[8]), .B(n8977), .Y(n1975) );
  INVX1 U8226 ( .A(n1975), .Y(n6820) );
  AND2X1 U8227 ( .A(recentdatapoints_head_i[24]), .B(n8979), .Y(n1959) );
  INVX1 U8228 ( .A(n1959), .Y(n6821) );
  AND2X1 U8229 ( .A(p_tmp_i_reg_1556[25]), .B(n8979), .Y(n1912) );
  INVX1 U8230 ( .A(n1912), .Y(n6822) );
  AND2X1 U8231 ( .A(p_tmp_i_reg_1556[13]), .B(n8980), .Y(n1888) );
  INVX1 U8232 ( .A(n1888), .Y(n6823) );
  AND2X1 U8233 ( .A(CircularBuffer_head_i_read_ass_reg_1624[10]), .B(n9011), 
        .Y(n1775) );
  INVX1 U8234 ( .A(n1775), .Y(n6824) );
  AND2X1 U8235 ( .A(recentVBools_head_i[14]), .B(n9010), .Y(n1762) );
  INVX1 U8236 ( .A(n1762), .Y(n6825) );
  AND2X1 U8237 ( .A(CircularBuffer_head_i_read_ass_reg_1624[22]), .B(n9009), 
        .Y(n1739) );
  INVX1 U8238 ( .A(n1739), .Y(n6826) );
  AND2X1 U8239 ( .A(CircularBuffer_head_i_read_ass_reg_1624[31]), .B(n9008), 
        .Y(n1712) );
  INVX1 U8240 ( .A(n1712), .Y(n6827) );
  AND2X1 U8241 ( .A(n2774), .B(n8991), .Y(n1633) );
  INVX1 U8242 ( .A(n1633), .Y(n6828) );
  BUFX2 U8243 ( .A(n2785), .Y(n6829) );
  BUFX2 U8244 ( .A(n2841), .Y(n6830) );
  BUFX2 U8245 ( .A(n2769), .Y(n6831) );
  BUFX2 U8246 ( .A(n2741), .Y(n6832) );
  AND2X1 U8247 ( .A(CircularBuffer_len_write_assig_fu_817_p2[4]), .B(n1646), 
        .Y(n1597) );
  INVX1 U8248 ( .A(n1597), .Y(n6833) );
  AND2X1 U8249 ( .A(CircularBuffer_len_write_assig_fu_817_p2[14]), .B(n8894), 
        .Y(n1581) );
  INVX1 U8250 ( .A(n1581), .Y(n6834) );
  AND2X1 U8251 ( .A(CircularBuffer_sum_read_assign_reg_1610[11]), .B(n9007), 
        .Y(n1444) );
  INVX1 U8252 ( .A(n1444), .Y(n6835) );
  AND2X1 U8253 ( .A(CircularBuffer_sum_read_assign_reg_1610[17]), .B(n9006), 
        .Y(n1432) );
  INVX1 U8254 ( .A(n1432), .Y(n6836) );
  AND2X1 U8255 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[10]), .Y(n2656) );
  INVX1 U8256 ( .A(n2656), .Y(n6837) );
  BUFX2 U8257 ( .A(n2721), .Y(n6838) );
  BUFX2 U8258 ( .A(n2709), .Y(n6839) );
  AND2X1 U8259 ( .A(n9012), .B(sum_phi_fu_311_p4[24]), .Y(n2600) );
  INVX1 U8260 ( .A(n2600), .Y(n6840) );
  AND2X1 U8261 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[16]), .B(n9040), 
        .Y(n1307) );
  INVX1 U8262 ( .A(n1307), .Y(n6841) );
  AND2X1 U8263 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[21]), .B(n9039), 
        .Y(n1295) );
  INVX1 U8264 ( .A(n1295), .Y(n6842) );
  AND2X1 U8265 ( .A(recentABools_head_i[26]), .B(n9038), .Y(n1281) );
  INVX1 U8266 ( .A(n1281), .Y(n6843) );
  AND2X1 U8267 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[31]), .B(n9037), 
        .Y(n1271) );
  INVX1 U8268 ( .A(n1271), .Y(n6844) );
  AND2X1 U8269 ( .A(tmp_5_fu_726_p2[4]), .B(n8992), .Y(n1192) );
  INVX1 U8270 ( .A(n1192), .Y(n6845) );
  AND2X1 U8271 ( .A(VbeatFallDelay_new_1_reg_342[7]), .B(n9013), .Y(n2164) );
  INVX1 U8272 ( .A(n2164), .Y(n6846) );
  AND2X1 U8273 ( .A(VbeatFallDelay[8]), .B(n9036), .Y(n1174) );
  INVX1 U8274 ( .A(n1174), .Y(n6847) );
  AND2X1 U8275 ( .A(tmp_5_fu_726_p2[11]), .B(n8993), .Y(n1164) );
  INVX1 U8276 ( .A(n1164), .Y(n6848) );
  AND2X1 U8277 ( .A(VbeatFallDelay[19]), .B(n9035), .Y(n1130) );
  INVX1 U8278 ( .A(n1130), .Y(n6849) );
  AND2X1 U8279 ( .A(VbeatFallDelay_new_1_reg_342[24]), .B(n9013), .Y(n2181) );
  INVX1 U8280 ( .A(n2181), .Y(n6850) );
  AND2X1 U8281 ( .A(tmp_5_fu_726_p2[29]), .B(n8994), .Y(n1092) );
  INVX1 U8282 ( .A(n1092), .Y(n6851) );
  AND2X1 U8283 ( .A(VbeatFallDelay[29]), .B(n9034), .Y(n1090) );
  INVX1 U8284 ( .A(n1090), .Y(n6852) );
  AND2X1 U8285 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[0]), .Y(n2566) );
  INVX1 U8286 ( .A(n2566), .Y(n6853) );
  AND2X1 U8287 ( .A(VbeatDelay[6]), .B(n9033), .Y(n1057) );
  INVX1 U8288 ( .A(n1057), .Y(n6854) );
  AND2X1 U8289 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[12]), .Y(n2554) );
  INVX1 U8290 ( .A(n2554), .Y(n6855) );
  AND2X1 U8291 ( .A(tmp_4_fu_716_p2[16]), .B(n8995), .Y(n1027) );
  INVX1 U8292 ( .A(n1027), .Y(n6856) );
  AND2X1 U8293 ( .A(VbeatDelay[18]), .B(n9032), .Y(n1017) );
  INVX1 U8294 ( .A(n1017), .Y(n6857) );
  AND2X1 U8295 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[24]), .Y(n2542) );
  INVX1 U8296 ( .A(n2542), .Y(n6858) );
  BUFX2 U8297 ( .A(n2332), .Y(n6859) );
  AND2X1 U8298 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[5]), .Y(n2426) );
  INVX1 U8299 ( .A(n2426), .Y(n6860) );
  AND2X1 U8300 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[14]), .Y(n2462) );
  INVX1 U8301 ( .A(n2462), .Y(n6861) );
  BUFX2 U8302 ( .A(n2318), .Y(n6862) );
  AND2X1 U8303 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[26]), .Y(n2510) );
  INVX1 U8304 ( .A(n2510), .Y(n6863) );
  BUFX2 U8305 ( .A(n2306), .Y(n6864) );
  AND2X1 U8306 ( .A(n2257), .B(n9019), .Y(n942) );
  INVX1 U8307 ( .A(n942), .Y(n6865) );
  BUFX2 U8308 ( .A(n2386), .Y(n6866) );
  BUFX2 U8309 ( .A(n2284), .Y(n6867) );
  BUFX2 U8310 ( .A(n2360), .Y(n6868) );
  AND2X1 U8311 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[4]), .B(n970), 
        .Y(n921) );
  INVX1 U8312 ( .A(n921), .Y(n6869) );
  AND2X1 U8313 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[14]), .B(n8891), .Y(n905) );
  INVX1 U8314 ( .A(n905), .Y(n6870) );
  AND2X1 U8315 ( .A(tmp_3_fu_706_p2[5]), .B(n8996), .Y(n775) );
  INVX1 U8316 ( .A(n775), .Y(n6871) );
  AND2X1 U8317 ( .A(AbeatDelay_new_reg_394[8]), .B(n9041), .Y(n2226) );
  INVX1 U8318 ( .A(n2226), .Y(n6872) );
  AND2X1 U8319 ( .A(AbeatDelay[17]), .B(n10670), .Y(n733) );
  INVX1 U8320 ( .A(n733), .Y(n6873) );
  AND2X1 U8321 ( .A(tmp_3_fu_706_p2[22]), .B(n8997), .Y(n719) );
  INVX1 U8322 ( .A(n719), .Y(n6874) );
  AND2X1 U8323 ( .A(AbeatDelay_new_reg_394[23]), .B(n9041), .Y(n2211) );
  INVX1 U8324 ( .A(n2211), .Y(n6875) );
  AND2X1 U8325 ( .A(AbeatDelay[30]), .B(n8896), .Y(n689) );
  INVX1 U8326 ( .A(n689), .Y(n6876) );
  AND2X1 U8327 ( .A(tmp_6_fu_497_p3[3]), .B(n8967), .Y(n675) );
  INVX1 U8328 ( .A(n675), .Y(n6877) );
  AND2X1 U8329 ( .A(AstimDelay[15]), .B(n8896), .Y(n638) );
  INVX1 U8330 ( .A(n638), .Y(n6878) );
  AND2X1 U8331 ( .A(tmp_6_fu_497_p3[17]), .B(n8966), .Y(n633) );
  INVX1 U8332 ( .A(n633), .Y(n6879) );
  AND2X1 U8333 ( .A(VstimDelay[1]), .B(n10670), .Y(n580) );
  INVX1 U8334 ( .A(n580), .Y(n6880) );
  AND2X1 U8335 ( .A(tmp_7_fu_511_p3[5]), .B(n8965), .Y(n569) );
  INVX1 U8336 ( .A(n569), .Y(n6881) );
  AND2X1 U8337 ( .A(tmp_7_fu_511_p3[21]), .B(n8964), .Y(n521) );
  INVX1 U8338 ( .A(n521), .Y(n6882) );
  AND2X1 U8339 ( .A(VstimDelay[24]), .B(n10670), .Y(n511) );
  INVX1 U8340 ( .A(n511), .Y(n6883) );
  AND2X1 U8341 ( .A(\Decision_AXILiteS_s_axi_U/n364 ), .B(
        \Decision_AXILiteS_s_axi_U/n351 ), .Y(\Decision_AXILiteS_s_axi_U/n363 ) );
  INVX1 U8342 ( .A(\Decision_AXILiteS_s_axi_U/n363 ), .Y(n6884) );
  AND2X1 U8343 ( .A(a_length[26]), .B(n8116), .Y(
        \Decision_AXILiteS_s_axi_U/n426 ) );
  INVX1 U8344 ( .A(\Decision_AXILiteS_s_axi_U/n426 ), .Y(n6885) );
  AND2X1 U8345 ( .A(\Decision_AXILiteS_s_axi_U/n368 ), .B(n8411), .Y(
        \Decision_AXILiteS_s_axi_U/n468 ) );
  INVX1 U8346 ( .A(\Decision_AXILiteS_s_axi_U/n468 ), .Y(n6886) );
  AND2X1 U8347 ( .A(\Decision_AXILiteS_s_axi_U/n356 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n514 ) );
  INVX1 U8348 ( .A(\Decision_AXILiteS_s_axi_U/n514 ), .Y(n6887) );
  AND2X1 U8349 ( .A(vthresh[27]), .B(n7865), .Y(
        \Decision_AXILiteS_s_axi_U/n488 ) );
  INVX1 U8350 ( .A(\Decision_AXILiteS_s_axi_U/n488 ), .Y(n6888) );
  AND2X1 U8351 ( .A(\Decision_AXILiteS_s_axi_U/n358 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n557 ) );
  INVX1 U8352 ( .A(\Decision_AXILiteS_s_axi_U/n557 ), .Y(n6889) );
  AND2X1 U8353 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[15]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n444 )
         );
  INVX1 U8354 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n444 ), 
        .Y(n6890) );
  AND2X1 U8355 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[14]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n476 )
         );
  INVX1 U8356 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n476 ), 
        .Y(n6891) );
  AND2X1 U8357 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[13]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n508 )
         );
  INVX1 U8358 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n508 ), 
        .Y(n6892) );
  AND2X1 U8359 ( .A(n9467), .B(data_read_reg_1495[12]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n540 )
         );
  INVX1 U8360 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n540 ), 
        .Y(n6893) );
  AND2X1 U8361 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][2] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n555 )
         );
  INVX1 U8362 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n555 ), 
        .Y(n6894) );
  AND2X1 U8363 ( .A(n9468), .B(data_read_reg_1495[5]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n594 )
         );
  INVX1 U8364 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n594 ), 
        .Y(n6895) );
  AND2X1 U8365 ( .A(n9468), .B(data_read_reg_1495[11]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n606 )
         );
  INVX1 U8366 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n606 ), 
        .Y(n6896) );
  AND2X1 U8367 ( .A(n9469), .B(data_read_reg_1495[4]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n626 )
         );
  INVX1 U8368 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n626 ), 
        .Y(n6897) );
  AND2X1 U8369 ( .A(n9469), .B(data_read_reg_1495[10]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n638 )
         );
  INVX1 U8370 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n638 ), 
        .Y(n6898) );
  AND2X1 U8371 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][15] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n705 )
         );
  INVX1 U8372 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n705 ), 
        .Y(n6899) );
  AND2X1 U8373 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][14] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n721 )
         );
  INVX1 U8374 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n721 ), 
        .Y(n6900) );
  AND2X1 U8375 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][1] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n725 )
         );
  INVX1 U8376 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n725 ), 
        .Y(n6901) );
  AND2X1 U8377 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][13] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n737 )
         );
  INVX1 U8378 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n737 ), 
        .Y(n6902) );
  AND2X1 U8379 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][0] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n741 )
         );
  INVX1 U8380 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n741 ), 
        .Y(n6903) );
  AND2X1 U8381 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][12] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n753 )
         );
  INVX1 U8382 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n753 ), 
        .Y(n6904) );
  AND2X1 U8383 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][11] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n769 )
         );
  INVX1 U8384 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n769 ), 
        .Y(n6905) );
  AND2X1 U8385 ( .A(n9466), .B(data_read_reg_1495[3]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n782 )
         );
  INVX1 U8386 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n782 ), 
        .Y(n6906) );
  AND2X1 U8387 ( .A(n9466), .B(data_read_reg_1495[9]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n794 )
         );
  INVX1 U8388 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n794 ), 
        .Y(n6907) );
  AND2X1 U8389 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][10] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n819 )
         );
  INVX1 U8390 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n819 ), 
        .Y(n6908) );
  AND2X1 U8391 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][9] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n836 )
         );
  INVX1 U8392 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n836 ), 
        .Y(n6909) );
  AND2X1 U8393 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][8] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n852 )
         );
  INVX1 U8394 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n852 ), 
        .Y(n6910) );
  AND2X1 U8395 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[2]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n866 )
         );
  INVX1 U8396 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n866 ), 
        .Y(n6911) );
  AND2X1 U8397 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[8]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n878 )
         );
  INVX1 U8398 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n878 ), 
        .Y(n6912) );
  AND2X1 U8399 ( .A(sum_1_reg_376[23]), .B(n8930), .Y(n2500) );
  INVX1 U8400 ( .A(n2500), .Y(n6913) );
  AND2X1 U8401 ( .A(sum_1_reg_376[0]), .B(n8930), .Y(n2408) );
  INVX1 U8402 ( .A(n2408), .Y(n6914) );
  AND2X1 U8403 ( .A(sum_reg_308[14]), .B(n8929), .Y(n2642) );
  INVX1 U8404 ( .A(n2642), .Y(n6915) );
  AND2X1 U8405 ( .A(sum_1_reg_376[9]), .B(n8930), .Y(n2444) );
  INVX1 U8406 ( .A(n2444), .Y(n6916) );
  AND2X1 U8407 ( .A(tmp_29_i_fu_752_p2[19]), .B(n8920), .Y(n3174) );
  INVX1 U8408 ( .A(n3174), .Y(n6917) );
  AND2X1 U8409 ( .A(tmp_29_i1_fu_1065_p2[19]), .B(n8922), .Y(n3226) );
  INVX1 U8410 ( .A(n3226), .Y(n6918) );
  AND2X1 U8411 ( .A(tmp_29_i_fu_752_p2[8]), .B(n8920), .Y(n3154) );
  INVX1 U8412 ( .A(n3154), .Y(n6919) );
  AND2X1 U8413 ( .A(tmp_29_i1_fu_1065_p2[8]), .B(n8922), .Y(n3206) );
  INVX1 U8414 ( .A(n3206), .Y(n6920) );
  AND2X1 U8415 ( .A(sum_reg_308[25]), .B(n8929), .Y(n2598) );
  INVX1 U8416 ( .A(n2598), .Y(n6921) );
  INVX1 U8417 ( .A(n4623), .Y(n6922) );
  AND2X1 U8418 ( .A(ACaptureThresh_loc_reg_288[11]), .B(n8969), .Y(n3040) );
  INVX1 U8419 ( .A(n3040), .Y(n6923) );
  BUFX2 U8420 ( .A(n3039), .Y(n6924) );
  INVX1 U8421 ( .A(n4607), .Y(n6925) );
  AND2X1 U8422 ( .A(ACaptureThresh_loc_reg_288[27]), .B(n8971), .Y(n3008) );
  INVX1 U8423 ( .A(n3008), .Y(n6926) );
  BUFX2 U8424 ( .A(n3007), .Y(n6927) );
  INVX1 U8425 ( .A(n4561), .Y(n6928) );
  AND2X1 U8426 ( .A(VCaptureThresh_loc_reg_298[9]), .B(n8970), .Y(n2916) );
  INVX1 U8427 ( .A(n2916), .Y(n6929) );
  BUFX2 U8428 ( .A(n2915), .Y(n6930) );
  INVX1 U8429 ( .A(n4546), .Y(n6931) );
  AND2X1 U8430 ( .A(VCaptureThresh_loc_reg_298[24]), .B(n8969), .Y(n2886) );
  INVX1 U8431 ( .A(n2886), .Y(n6932) );
  BUFX2 U8432 ( .A(n2885), .Y(n6933) );
  BUFX2 U8433 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n29 ), 
        .Y(n6934) );
  BUFX2 U8434 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n30 ), 
        .Y(n6935) );
  AND2X1 U8435 ( .A(n9939), .B(n9938), .Y(n1820) );
  INVX1 U8436 ( .A(n1820), .Y(n6936) );
  AND2X1 U8437 ( .A(n10247), .B(n10246), .Y(n1264) );
  INVX1 U8438 ( .A(n1264), .Y(n6937) );
  AND2X1 U8439 ( .A(n10527), .B(n10457), .Y(n339) );
  INVX1 U8440 ( .A(n339), .Y(n6938) );
  AND2X1 U8441 ( .A(n9844), .B(n9845), .Y(n2038) );
  INVX1 U8442 ( .A(n2038), .Y(n6939) );
  AND2X1 U8443 ( .A(n9870), .B(n9869), .Y(n1941) );
  INVX1 U8444 ( .A(n1941), .Y(n6940) );
  AND2X1 U8445 ( .A(recentdatapoints_len_load_op_fu_556_p2[6]), .B(n8972), .Y(
        n1826) );
  INVX1 U8446 ( .A(n1826), .Y(n6941) );
  AND2X1 U8447 ( .A(recentdatapoints_len_load_op_fu_556_p2[20]), .B(n8972), 
        .Y(n1843) );
  INVX1 U8448 ( .A(n1843), .Y(n6942) );
  AND2X1 U8449 ( .A(n9886), .B(n8976), .Y(n1861) );
  INVX1 U8450 ( .A(n1861), .Y(n6943) );
  AND2X1 U8451 ( .A(recentdatapoints_data_q0[1]), .B(n8869), .Y(n416) );
  INVX1 U8452 ( .A(n416), .Y(n6944) );
  AND2X1 U8453 ( .A(recentdatapoints_data_q0[14]), .B(n8868), .Y(n419) );
  INVX1 U8454 ( .A(n419), .Y(n6945) );
  AND2X1 U8455 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[3]), 
        .Y(n454) );
  INVX1 U8456 ( .A(n454), .Y(n6946) );
  AND2X1 U8457 ( .A(CircularBuffer_len_read_assign_fu_772_p2[25]), .B(n8919), 
        .Y(n2744) );
  INVX1 U8458 ( .A(n2744), .Y(n6947) );
  AND2X1 U8459 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[25]), .B(n8921), .Y(n2251) );
  INVX1 U8460 ( .A(n2251), .Y(n6948) );
  AND2X1 U8461 ( .A(n8881), .B(\Decision_AXILiteS_s_axi_U/n396 ), .Y(
        \Decision_AXILiteS_s_axi_U/n388 ) );
  INVX1 U8462 ( .A(\Decision_AXILiteS_s_axi_U/n388 ), .Y(n6949) );
  AND2X1 U8463 ( .A(\Decision_AXILiteS_s_axi_U/n429 ), .B(
        \Decision_AXILiteS_s_axi_U/n352 ), .Y(\Decision_AXILiteS_s_axi_U/n442 ) );
  INVX1 U8464 ( .A(\Decision_AXILiteS_s_axi_U/n442 ), .Y(n6950) );
  OR2X1 U8465 ( .A(AbeatDelay_new_reg_394[13]), .B(AbeatDelay_new_reg_394[12]), 
        .Y(n11057) );
  INVX1 U8466 ( .A(n11057), .Y(n6951) );
  OR2X1 U8467 ( .A(AbeatDelay_new_reg_394[15]), .B(AbeatDelay_new_reg_394[14]), 
        .Y(n11056) );
  INVX1 U8468 ( .A(n11056), .Y(n6952) );
  AND2X1 U8469 ( .A(v_flip[6]), .B(n8951), .Y(n3128) );
  INVX1 U8470 ( .A(n3128), .Y(n6953) );
  AND2X1 U8471 ( .A(a_length[6]), .B(n8952), .Y(n3114) );
  INVX1 U8472 ( .A(n3114), .Y(n6954) );
  AND2X1 U8473 ( .A(a_length[26]), .B(n8953), .Y(n3074) );
  INVX1 U8474 ( .A(n3074), .Y(n6955) );
  AND2X1 U8475 ( .A(v_length[18]), .B(n8955), .Y(n2962) );
  INVX1 U8476 ( .A(n2962), .Y(n6956) );
  AND2X1 U8477 ( .A(v_length[28]), .B(n8954), .Y(n2942) );
  INVX1 U8478 ( .A(n2942), .Y(n6957) );
  AND2X1 U8479 ( .A(recentdatapoints_head_i[14]), .B(n8980), .Y(n1969) );
  INVX1 U8480 ( .A(n1969), .Y(n6958) );
  AND2X1 U8481 ( .A(recentdatapoints_head_i[25]), .B(n8980), .Y(n1958) );
  INVX1 U8482 ( .A(n1958), .Y(n6959) );
  AND2X1 U8483 ( .A(n8963), .B(recentdatapoints_head_i[4]), .Y(n1930) );
  INVX1 U8484 ( .A(n1930), .Y(n6960) );
  AND2X1 U8485 ( .A(p_tmp_i_reg_1556[24]), .B(n8979), .Y(n1910) );
  INVX1 U8486 ( .A(n1910), .Y(n6961) );
  AND2X1 U8487 ( .A(p_tmp_i_reg_1556[11]), .B(n8978), .Y(n1884) );
  INVX1 U8488 ( .A(n1884), .Y(n6962) );
  AND2X1 U8489 ( .A(recentVBools_head_i[10]), .B(n9011), .Y(n1774) );
  INVX1 U8490 ( .A(n1774), .Y(n6963) );
  AND2X1 U8491 ( .A(CircularBuffer_head_i_read_ass_reg_1624[15]), .B(n9010), 
        .Y(n1760) );
  INVX1 U8492 ( .A(n1760), .Y(n6964) );
  AND2X1 U8493 ( .A(CircularBuffer_head_i_read_ass_reg_1624[24]), .B(n9009), 
        .Y(n1733) );
  INVX1 U8494 ( .A(n1733), .Y(n6965) );
  AND2X1 U8495 ( .A(recentVBools_head_i[31]), .B(n9008), .Y(n1711) );
  INVX1 U8496 ( .A(n1711), .Y(n6966) );
  AND2X1 U8497 ( .A(n2766), .B(n8992), .Y(n1627) );
  INVX1 U8498 ( .A(n1627), .Y(n6967) );
  BUFX2 U8499 ( .A(n2783), .Y(n6968) );
  BUFX2 U8500 ( .A(n2839), .Y(n6969) );
  BUFX2 U8501 ( .A(n2767), .Y(n6970) );
  BUFX2 U8502 ( .A(n2823), .Y(n6971) );
  AND2X1 U8503 ( .A(CircularBuffer_len_write_assig_fu_817_p2[5]), .B(n1646), 
        .Y(n1596) );
  INVX1 U8504 ( .A(n1596), .Y(n6972) );
  AND2X1 U8505 ( .A(CircularBuffer_len_write_assig_fu_817_p2[15]), .B(n8894), 
        .Y(n1580) );
  INVX1 U8506 ( .A(n1580), .Y(n6973) );
  AND2X1 U8507 ( .A(CircularBuffer_sum_read_assign_reg_1610[16]), .B(n9007), 
        .Y(n1434) );
  INVX1 U8508 ( .A(n1434), .Y(n6974) );
  AND2X1 U8509 ( .A(CircularBuffer_sum_read_assign_reg_1610[20]), .B(n9006), 
        .Y(n1426) );
  INVX1 U8510 ( .A(n1426), .Y(n6975) );
  BUFX2 U8511 ( .A(n2733), .Y(n6976) );
  AND2X1 U8512 ( .A(n9012), .B(sum_phi_fu_311_p4[11]), .Y(n2652) );
  INVX1 U8513 ( .A(n2652), .Y(n6977) );
  BUFX2 U8514 ( .A(n2720), .Y(n6978) );
  AND2X1 U8515 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[25]), .Y(n2596) );
  INVX1 U8516 ( .A(n2596), .Y(n6979) );
  BUFX2 U8517 ( .A(n2707), .Y(n6980) );
  AND2X1 U8518 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[11]), .B(n9034), 
        .Y(n1362) );
  INVX1 U8519 ( .A(n1362), .Y(n6981) );
  AND2X1 U8520 ( .A(recentABools_head_i[0]), .B(ap_CS_fsm[7]), .Y(n1336) );
  INVX1 U8521 ( .A(n1336), .Y(n6982) );
  AND2X1 U8522 ( .A(recentABools_head_i[16]), .B(n9040), .Y(n1306) );
  INVX1 U8523 ( .A(n1306), .Y(n6983) );
  AND2X1 U8524 ( .A(recentABools_head_i[21]), .B(n9039), .Y(n1294) );
  INVX1 U8525 ( .A(n1294), .Y(n6984) );
  AND2X1 U8526 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[27]), .B(n9038), 
        .Y(n1279) );
  INVX1 U8527 ( .A(n1279), .Y(n6985) );
  AND2X1 U8528 ( .A(VbeatFallDelay[3]), .B(n9037), .Y(n1194) );
  INVX1 U8529 ( .A(n1194), .Y(n6986) );
  AND2X1 U8530 ( .A(VbeatFallDelay_new_1_reg_342[9]), .B(n9013), .Y(n2166) );
  INVX1 U8531 ( .A(n2166), .Y(n6987) );
  AND2X1 U8532 ( .A(VbeatFallDelay[11]), .B(n9036), .Y(n1162) );
  INVX1 U8533 ( .A(n1162), .Y(n6988) );
  AND2X1 U8534 ( .A(tmp_5_fu_726_p2[12]), .B(n8993), .Y(n1160) );
  INVX1 U8535 ( .A(n1160), .Y(n6989) );
  AND2X1 U8536 ( .A(VbeatFallDelay_new_1_reg_342[25]), .B(n9013), .Y(n2182) );
  INVX1 U8537 ( .A(n2182), .Y(n6990) );
  AND2X1 U8538 ( .A(tmp_5_fu_726_p2[30]), .B(n8994), .Y(n1088) );
  INVX1 U8539 ( .A(n1088), .Y(n6991) );
  AND2X1 U8540 ( .A(VbeatDelay[0]), .B(n9033), .Y(n1076) );
  INVX1 U8541 ( .A(n1076), .Y(n6992) );
  AND2X1 U8542 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[1]), .Y(n2565) );
  INVX1 U8543 ( .A(n2565), .Y(n6993) );
  AND2X1 U8544 ( .A(VbeatDelay[11]), .B(n9032), .Y(n1041) );
  INVX1 U8545 ( .A(n1041), .Y(n6994) );
  AND2X1 U8546 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[13]), .Y(n2553) );
  INVX1 U8547 ( .A(n2553), .Y(n6995) );
  AND2X1 U8548 ( .A(tmp_4_fu_716_p2[17]), .B(n8995), .Y(n1023) );
  INVX1 U8549 ( .A(n1023), .Y(n6996) );
  AND2X1 U8550 ( .A(VbeatDelay[20]), .B(n9035), .Y(n1011) );
  INVX1 U8551 ( .A(n1011), .Y(n6997) );
  AND2X1 U8552 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[25]), .Y(n2541) );
  INVX1 U8553 ( .A(n2541), .Y(n6998) );
  AND2X1 U8554 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[6]), .Y(n2430) );
  INVX1 U8555 ( .A(n2430), .Y(n6999) );
  BUFX2 U8556 ( .A(n2324), .Y(n7000) );
  AND2X1 U8557 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[16]), .Y(n2470) );
  INVX1 U8558 ( .A(n2470), .Y(n7001) );
  BUFX2 U8559 ( .A(n2309), .Y(n7002) );
  AND2X1 U8560 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[27]), .Y(n2514) );
  INVX1 U8561 ( .A(n2514), .Y(n7003) );
  AND2X1 U8562 ( .A(n9017), .B(CircularBuffer_len_read_assign_3_fu_1091_p3[1]), 
        .Y(n968) );
  INVX1 U8563 ( .A(n968), .Y(n7004) );
  AND2X1 U8564 ( .A(n2279), .B(n9019), .Y(n955) );
  INVX1 U8565 ( .A(n955), .Y(n7005) );
  BUFX2 U8566 ( .A(n2296), .Y(n7006) );
  BUFX2 U8567 ( .A(n2384), .Y(n7007) );
  BUFX2 U8568 ( .A(n2274), .Y(n7008) );
  BUFX2 U8569 ( .A(n2358), .Y(n7009) );
  AND2X1 U8570 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[5]), .B(n970), 
        .Y(n920) );
  INVX1 U8571 ( .A(n920), .Y(n7010) );
  AND2X1 U8572 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[15]), .B(n8891), .Y(n904) );
  INVX1 U8573 ( .A(n904), .Y(n7011) );
  AND2X1 U8574 ( .A(tmp_3_fu_706_p2[6]), .B(n8996), .Y(n772) );
  INVX1 U8575 ( .A(n772), .Y(n7012) );
  AND2X1 U8576 ( .A(AbeatDelay_new_reg_394[10]), .B(n9041), .Y(n2224) );
  INVX1 U8577 ( .A(n2224), .Y(n7013) );
  AND2X1 U8578 ( .A(AbeatDelay[11]), .B(n8896), .Y(n755) );
  INVX1 U8579 ( .A(n755), .Y(n7014) );
  AND2X1 U8580 ( .A(AbeatDelay_new_reg_394[24]), .B(n9041), .Y(n2210) );
  INVX1 U8581 ( .A(n2210), .Y(n7015) );
  AND2X1 U8582 ( .A(tmp_3_fu_706_p2[25]), .B(n8997), .Y(n708) );
  INVX1 U8583 ( .A(n708), .Y(n7016) );
  AND2X1 U8584 ( .A(AbeatDelay[31]), .B(n8896), .Y(n686) );
  INVX1 U8585 ( .A(n686), .Y(n7017) );
  AND2X1 U8586 ( .A(tmp_6_fu_497_p3[4]), .B(n8967), .Y(n672) );
  INVX1 U8587 ( .A(n672), .Y(n7018) );
  AND2X1 U8588 ( .A(AstimDelay[16]), .B(n8896), .Y(n635) );
  INVX1 U8589 ( .A(n635), .Y(n7019) );
  AND2X1 U8590 ( .A(tmp_6_fu_497_p3[20]), .B(n8966), .Y(n624) );
  INVX1 U8591 ( .A(n624), .Y(n7020) );
  AND2X1 U8592 ( .A(VstimDelay[2]), .B(n8896), .Y(n577) );
  INVX1 U8593 ( .A(n577), .Y(n7021) );
  AND2X1 U8594 ( .A(tmp_7_fu_511_p3[6]), .B(n8965), .Y(n566) );
  INVX1 U8595 ( .A(n566), .Y(n7022) );
  AND2X1 U8596 ( .A(tmp_7_fu_511_p3[22]), .B(n8964), .Y(n518) );
  INVX1 U8597 ( .A(n518), .Y(n7023) );
  AND2X1 U8598 ( .A(VstimDelay[25]), .B(n8896), .Y(n508) );
  INVX1 U8599 ( .A(n508), .Y(n7024) );
  AND2X1 U8600 ( .A(a_length[29]), .B(n8116), .Y(
        \Decision_AXILiteS_s_axi_U/n423 ) );
  INVX1 U8601 ( .A(\Decision_AXILiteS_s_axi_U/n423 ), .Y(n7025) );
  AND2X1 U8602 ( .A(\Decision_AXILiteS_s_axi_U/n366 ), .B(n8411), .Y(
        \Decision_AXILiteS_s_axi_U/n467 ) );
  INVX1 U8603 ( .A(\Decision_AXILiteS_s_axi_U/n467 ), .Y(n7026) );
  AND2X1 U8604 ( .A(\Decision_AXILiteS_s_axi_U/n358 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n515 ) );
  INVX1 U8605 ( .A(\Decision_AXILiteS_s_axi_U/n515 ), .Y(n7027) );
  AND2X1 U8606 ( .A(vthresh[28]), .B(n7865), .Y(
        \Decision_AXILiteS_s_axi_U/n487 ) );
  INVX1 U8607 ( .A(\Decision_AXILiteS_s_axi_U/n487 ), .Y(n7028) );
  AND2X1 U8608 ( .A(\Decision_AXILiteS_s_axi_U/n356 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n556 ) );
  INVX1 U8609 ( .A(\Decision_AXILiteS_s_axi_U/n556 ), .Y(n7029) );
  AND2X1 U8610 ( .A(s_axi_AXILiteS_AWADDR[0]), .B(n8652), .Y(
        \Decision_AXILiteS_s_axi_U/n635 ) );
  INVX1 U8611 ( .A(\Decision_AXILiteS_s_axi_U/n635 ), .Y(n7030) );
  AND2X1 U8612 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[14]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n442 )
         );
  INVX1 U8613 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n442 ), 
        .Y(n7031) );
  AND2X1 U8614 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[15]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n478 )
         );
  INVX1 U8615 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n478 ), 
        .Y(n7032) );
  AND2X1 U8616 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[12]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n506 )
         );
  INVX1 U8617 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n506 ), 
        .Y(n7033) );
  AND2X1 U8618 ( .A(n9467), .B(data_read_reg_1495[13]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n542 )
         );
  INVX1 U8619 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n542 ), 
        .Y(n7034) );
  AND2X1 U8620 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][3] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n557 )
         );
  INVX1 U8621 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n557 ), 
        .Y(n7035) );
  AND2X1 U8622 ( .A(n9468), .B(data_read_reg_1495[4]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n592 )
         );
  INVX1 U8623 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n592 ), 
        .Y(n7036) );
  AND2X1 U8624 ( .A(n9468), .B(data_read_reg_1495[10]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n604 )
         );
  INVX1 U8625 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n604 ), 
        .Y(n7037) );
  AND2X1 U8626 ( .A(n9469), .B(data_read_reg_1495[5]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n628 )
         );
  INVX1 U8627 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n628 ), 
        .Y(n7038) );
  AND2X1 U8628 ( .A(n9469), .B(data_read_reg_1495[11]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n640 )
         );
  INVX1 U8629 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n640 ), 
        .Y(n7039) );
  AND2X1 U8630 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][14] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n704 )
         );
  INVX1 U8631 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n704 ), 
        .Y(n7040) );
  AND2X1 U8632 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][15] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n722 )
         );
  INVX1 U8633 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n722 ), 
        .Y(n7041) );
  AND2X1 U8634 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][0] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n724 )
         );
  INVX1 U8635 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n724 ), 
        .Y(n7042) );
  AND2X1 U8636 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][12] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n736 )
         );
  INVX1 U8637 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n736 ), 
        .Y(n7043) );
  AND2X1 U8638 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][1] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n742 )
         );
  INVX1 U8639 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n742 ), 
        .Y(n7044) );
  AND2X1 U8640 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][13] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n754 )
         );
  INVX1 U8641 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n754 ), 
        .Y(n7045) );
  AND2X1 U8642 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][10] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n768 )
         );
  INVX1 U8643 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n768 ), 
        .Y(n7046) );
  AND2X1 U8644 ( .A(n9466), .B(data_read_reg_1495[2]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n780 )
         );
  INVX1 U8645 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n780 ), 
        .Y(n7047) );
  AND2X1 U8646 ( .A(n9466), .B(data_read_reg_1495[8]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n792 )
         );
  INVX1 U8647 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n792 ), 
        .Y(n7048) );
  AND2X1 U8648 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][11] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n820 )
         );
  INVX1 U8649 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n820 ), 
        .Y(n7049) );
  AND2X1 U8650 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][8] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n835 )
         );
  INVX1 U8651 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n835 ), 
        .Y(n7050) );
  AND2X1 U8652 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][9] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n853 )
         );
  INVX1 U8653 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n853 ), 
        .Y(n7051) );
  AND2X1 U8654 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[3]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n868 )
         );
  INVX1 U8655 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n868 ), 
        .Y(n7052) );
  AND2X1 U8656 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[9]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n880 )
         );
  INVX1 U8657 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n880 ), 
        .Y(n7053) );
  BUFX2 U8658 ( .A(n12100), .Y(n7054) );
  AND2X1 U8659 ( .A(v_thresh[20]), .B(n9540), .Y(n12238) );
  INVX1 U8660 ( .A(n12238), .Y(n7055) );
  AND2X1 U8661 ( .A(a_thresh[20]), .B(n9490), .Y(n11605) );
  INVX1 U8662 ( .A(n11605), .Y(n7056) );
  AND2X1 U8663 ( .A(sum_reg_308[10]), .B(n8929), .Y(n2658) );
  INVX1 U8664 ( .A(n2658), .Y(n7057) );
  AND2X1 U8665 ( .A(sum_1_reg_376[30]), .B(n8930), .Y(n2528) );
  INVX1 U8666 ( .A(n2528), .Y(n7058) );
  AND2X1 U8667 ( .A(tmp_29_i_fu_752_p2[18]), .B(n8920), .Y(n3175) );
  INVX1 U8668 ( .A(n3175), .Y(n7059) );
  AND2X1 U8669 ( .A(tmp_29_i1_fu_1065_p2[18]), .B(n8922), .Y(n3227) );
  INVX1 U8670 ( .A(n3227), .Y(n7060) );
  AND2X1 U8671 ( .A(tmp_29_i_fu_752_p2[7]), .B(n8920), .Y(n3155) );
  INVX1 U8672 ( .A(n3155), .Y(n7061) );
  AND2X1 U8673 ( .A(tmp_29_i1_fu_1065_p2[7]), .B(n8922), .Y(n3207) );
  INVX1 U8674 ( .A(n3207), .Y(n7062) );
  AND2X1 U8675 ( .A(sum_1_reg_376[14]), .B(n8930), .Y(n2464) );
  INVX1 U8676 ( .A(n2464), .Y(n7063) );
  AND2X1 U8677 ( .A(sum_reg_308[22]), .B(n8929), .Y(n2610) );
  INVX1 U8678 ( .A(n2610), .Y(n7064) );
  INVX1 U8679 ( .A(n4621), .Y(n7065) );
  AND2X1 U8680 ( .A(ACaptureThresh_loc_reg_288[13]), .B(n8970), .Y(n3036) );
  INVX1 U8681 ( .A(n3036), .Y(n7066) );
  BUFX2 U8682 ( .A(n3035), .Y(n7067) );
  INVX1 U8683 ( .A(n4606), .Y(n7068) );
  AND2X1 U8684 ( .A(ACaptureThresh_loc_reg_288[28]), .B(n8971), .Y(n3006) );
  INVX1 U8685 ( .A(n3006), .Y(n7069) );
  BUFX2 U8686 ( .A(n3005), .Y(n7070) );
  INVX1 U8687 ( .A(n4560), .Y(n7071) );
  AND2X1 U8688 ( .A(VCaptureThresh_loc_reg_298[10]), .B(n8970), .Y(n2914) );
  INVX1 U8689 ( .A(n2914), .Y(n7072) );
  BUFX2 U8690 ( .A(n2913), .Y(n7073) );
  INVX1 U8691 ( .A(n4545), .Y(n7074) );
  AND2X1 U8692 ( .A(VCaptureThresh_loc_reg_298[25]), .B(n8969), .Y(n2884) );
  INVX1 U8693 ( .A(n2884), .Y(n7075) );
  BUFX2 U8694 ( .A(n2883), .Y(n7076) );
  AND2X1 U8695 ( .A(\toReturn_5_reg_1655[0] ), .B(n10057), .Y(n1469) );
  INVX1 U8696 ( .A(n1469), .Y(n7077) );
  BUFX2 U8697 ( .A(n1471), .Y(n7078) );
  AND2X1 U8698 ( .A(\toReturn_7_reg_1750[0] ), .B(n10535), .Y(n834) );
  INVX1 U8699 ( .A(n834), .Y(n7079) );
  BUFX2 U8700 ( .A(n836), .Y(n7080) );
  BUFX2 U8701 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n24 ), 
        .Y(n7081) );
  BUFX2 U8702 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n25 ), 
        .Y(n7082) );
  BUFX2 U8703 ( .A(\Decision_AXILiteS_s_axi_U/n370 ), .Y(n7083) );
  OR2X1 U8704 ( .A(n10899), .B(n10898), .Y(\Decision_AXILiteS_s_axi_U/n372 )
         );
  INVX1 U8705 ( .A(\Decision_AXILiteS_s_axi_U/n372 ), .Y(n7084) );
  BUFX2 U8706 ( .A(n278), .Y(n7085) );
  AND2X1 U8707 ( .A(n9873), .B(n9872), .Y(n1942) );
  INVX1 U8708 ( .A(n1942), .Y(n7086) );
  AND2X1 U8709 ( .A(n9955), .B(n9954), .Y(n1810) );
  INVX1 U8710 ( .A(n1810), .Y(n7087) );
  AND2X1 U8711 ( .A(n10263), .B(n10262), .Y(n1246) );
  INVX1 U8712 ( .A(n1246), .Y(n7088) );
  AND2X1 U8713 ( .A(n10499), .B(n10501), .Y(n322) );
  INVX1 U8714 ( .A(n322), .Y(n7089) );
  AND2X1 U8715 ( .A(n9847), .B(n9848), .Y(n2037) );
  INVX1 U8716 ( .A(n2037), .Y(n7090) );
  AND2X1 U8717 ( .A(recentdatapoints_len_load_op_fu_556_p2[7]), .B(n8972), .Y(
        n1827) );
  INVX1 U8718 ( .A(n1827), .Y(n7091) );
  AND2X1 U8719 ( .A(recentdatapoints_len_load_op_fu_556_p2[21]), .B(n8972), 
        .Y(n1845) );
  INVX1 U8720 ( .A(n1845), .Y(n7092) );
  AND2X1 U8721 ( .A(p_tmp_i_fu_587_p3[1]), .B(n8975), .Y(n1863) );
  INVX1 U8722 ( .A(n1863), .Y(n7093) );
  AND2X1 U8723 ( .A(CircularBuffer_len_read_assign_fu_772_p2[31]), .B(n3151), 
        .Y(n2862) );
  INVX1 U8724 ( .A(n2862), .Y(n7094) );
  AND2X1 U8725 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[31]), .B(n3149), .Y(n2401) );
  INVX1 U8726 ( .A(n2401), .Y(n7095) );
  AND2X1 U8727 ( .A(recentdatapoints_data_q0[7]), .B(n8869), .Y(n404) );
  INVX1 U8728 ( .A(n404), .Y(n7096) );
  AND2X1 U8729 ( .A(recentdatapoints_data_q0[10]), .B(n8868), .Y(n427) );
  INVX1 U8730 ( .A(n427), .Y(n7097) );
  AND2X1 U8731 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[13]), 
        .Y(n463) );
  INVX1 U8732 ( .A(n463), .Y(n7098) );
  AND2X1 U8733 ( .A(CircularBuffer_len_read_assign_fu_772_p2[22]), .B(n8919), 
        .Y(n2750) );
  INVX1 U8734 ( .A(n2750), .Y(n7099) );
  AND2X1 U8735 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[22]), .B(n8921), .Y(n2257) );
  INVX1 U8736 ( .A(n2257), .Y(n7100) );
  AND2X1 U8737 ( .A(n4695), .B(\tmp_s_reg_1578[0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n75 ) );
  INVX1 U8738 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n75 ), 
        .Y(n7101) );
  AND2X1 U8739 ( .A(n8881), .B(\Decision_AXILiteS_s_axi_U/n352 ), .Y(
        \Decision_AXILiteS_s_axi_U/n400 ) );
  INVX1 U8740 ( .A(\Decision_AXILiteS_s_axi_U/n400 ), .Y(n7102) );
  AND2X1 U8741 ( .A(\Decision_AXILiteS_s_axi_U/n429 ), .B(
        \Decision_AXILiteS_s_axi_U/n396 ), .Y(\Decision_AXILiteS_s_axi_U/n432 ) );
  INVX1 U8742 ( .A(\Decision_AXILiteS_s_axi_U/n432 ), .Y(n7103) );
  AND2X1 U8743 ( .A(v_flip[7]), .B(n8951), .Y(n3127) );
  INVX1 U8744 ( .A(n3127), .Y(n7104) );
  AND2X1 U8745 ( .A(a_length[5]), .B(n8952), .Y(n3116) );
  INVX1 U8746 ( .A(n3116), .Y(n7105) );
  AND2X1 U8747 ( .A(a_length[27]), .B(n8953), .Y(n3072) );
  INVX1 U8748 ( .A(n3072), .Y(n7106) );
  AND2X1 U8749 ( .A(v_length[19]), .B(n8955), .Y(n2960) );
  INVX1 U8750 ( .A(n2960), .Y(n7107) );
  AND2X1 U8751 ( .A(v_length[29]), .B(n8954), .Y(n2940) );
  INVX1 U8752 ( .A(n2940), .Y(n7108) );
  AND2X1 U8753 ( .A(recentdatapoints_head_i[15]), .B(n8980), .Y(n1968) );
  INVX1 U8754 ( .A(n1968), .Y(n7109) );
  AND2X1 U8755 ( .A(recentdatapoints_head_i[26]), .B(n8977), .Y(n1957) );
  INVX1 U8756 ( .A(n1957), .Y(n7110) );
  AND2X1 U8757 ( .A(p_tmp_i_reg_1556[23]), .B(n8979), .Y(n1908) );
  INVX1 U8758 ( .A(n1908), .Y(n7111) );
  AND2X1 U8759 ( .A(p_tmp_i_reg_1556[10]), .B(n8978), .Y(n1882) );
  INVX1 U8760 ( .A(n1882), .Y(n7112) );
  AND2X1 U8761 ( .A(CircularBuffer_head_i_read_ass_reg_1624[11]), .B(n9011), 
        .Y(n1772) );
  INVX1 U8762 ( .A(n1772), .Y(n7113) );
  AND2X1 U8763 ( .A(recentVBools_head_i[17]), .B(n9010), .Y(n1753) );
  INVX1 U8764 ( .A(n1753), .Y(n7114) );
  AND2X1 U8765 ( .A(recentVBools_head_i[22]), .B(n9009), .Y(n1738) );
  INVX1 U8766 ( .A(n1738), .Y(n7115) );
  AND2X1 U8767 ( .A(recentVBools_head_i[28]), .B(n9008), .Y(n1720) );
  INVX1 U8768 ( .A(n1720), .Y(n7116) );
  AND2X1 U8769 ( .A(n8991), .B(CircularBuffer_len_read_assign_1_fu_778_p3[4]), 
        .Y(n1641) );
  INVX1 U8770 ( .A(n1641), .Y(n7117) );
  AND2X1 U8771 ( .A(n2770), .B(n8992), .Y(n1630) );
  INVX1 U8772 ( .A(n1630), .Y(n7118) );
  BUFX2 U8773 ( .A(n2777), .Y(n7119) );
  BUFX2 U8774 ( .A(n2837), .Y(n7120) );
  BUFX2 U8775 ( .A(n2759), .Y(n7121) );
  BUFX2 U8776 ( .A(n2819), .Y(n7122) );
  AND2X1 U8777 ( .A(CircularBuffer_sum_read_assign_reg_1610[12]), .B(n9007), 
        .Y(n1442) );
  INVX1 U8778 ( .A(n1442), .Y(n7123) );
  AND2X1 U8779 ( .A(CircularBuffer_sum_read_assign_reg_1610[21]), .B(n9006), 
        .Y(n1424) );
  INVX1 U8780 ( .A(n1424), .Y(n7124) );
  BUFX2 U8781 ( .A(n2732), .Y(n7125) );
  AND2X1 U8782 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[12]), .Y(n2648) );
  INVX1 U8783 ( .A(n2648), .Y(n7126) );
  BUFX2 U8784 ( .A(n2718), .Y(n7127) );
  BUFX2 U8785 ( .A(n2706), .Y(n7128) );
  AND2X1 U8786 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[27]), .Y(n2588) );
  INVX1 U8787 ( .A(n2588), .Y(n7129) );
  AND2X1 U8788 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[25]), .B(n9031), 
        .Y(n1390) );
  INVX1 U8789 ( .A(n1390), .Y(n7130) );
  AND2X1 U8790 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[0]), .B(n9037), 
        .Y(n1340) );
  INVX1 U8791 ( .A(n1340), .Y(n7131) );
  AND2X1 U8792 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[17]), .B(n9040), 
        .Y(n1305) );
  INVX1 U8793 ( .A(n1305), .Y(n7132) );
  AND2X1 U8794 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[22]), .B(n9039), 
        .Y(n1292) );
  INVX1 U8795 ( .A(n1292), .Y(n7133) );
  AND2X1 U8796 ( .A(recentABools_head_i[27]), .B(n9038), .Y(n1278) );
  INVX1 U8797 ( .A(n1278), .Y(n7134) );
  AND2X1 U8798 ( .A(VbeatFallDelay[9]), .B(n9036), .Y(n1170) );
  INVX1 U8799 ( .A(n1170), .Y(n7135) );
  AND2X1 U8800 ( .A(VbeatFallDelay_new_1_reg_342[12]), .B(n9013), .Y(n2169) );
  INVX1 U8801 ( .A(n2169), .Y(n7136) );
  AND2X1 U8802 ( .A(tmp_5_fu_726_p2[13]), .B(n8993), .Y(n1156) );
  INVX1 U8803 ( .A(n1156), .Y(n7137) );
  AND2X1 U8804 ( .A(VbeatFallDelay[20]), .B(n9035), .Y(n1126) );
  INVX1 U8805 ( .A(n1126), .Y(n7138) );
  AND2X1 U8806 ( .A(VbeatFallDelay_new_1_reg_342[26]), .B(n9013), .Y(n2183) );
  INVX1 U8807 ( .A(n2183), .Y(n7139) );
  AND2X1 U8808 ( .A(VbeatFallDelay[30]), .B(n9034), .Y(n1086) );
  INVX1 U8809 ( .A(n1086), .Y(n7140) );
  AND2X1 U8810 ( .A(tmp_5_fu_726_p2[31]), .B(n8994), .Y(n1084) );
  INVX1 U8811 ( .A(n1084), .Y(n7141) );
  AND2X1 U8812 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[2]), .Y(n2564) );
  INVX1 U8813 ( .A(n2564), .Y(n7142) );
  AND2X1 U8814 ( .A(VbeatDelay[9]), .B(n9032), .Y(n1048) );
  INVX1 U8815 ( .A(n1048), .Y(n7143) );
  AND2X1 U8816 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[16]), .Y(n2550) );
  INVX1 U8817 ( .A(n2550), .Y(n7144) );
  AND2X1 U8818 ( .A(tmp_4_fu_716_p2[18]), .B(n8995), .Y(n1019) );
  INVX1 U8819 ( .A(n1019), .Y(n7145) );
  AND2X1 U8820 ( .A(VbeatDelay[19]), .B(n9033), .Y(n1014) );
  INVX1 U8821 ( .A(n1014), .Y(n7146) );
  AND2X1 U8822 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[26]), .Y(n2540) );
  INVX1 U8823 ( .A(n2540), .Y(n7147) );
  BUFX2 U8824 ( .A(n2331), .Y(n7148) );
  BUFX2 U8825 ( .A(n2319), .Y(n7149) );
  AND2X1 U8826 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[15]), .Y(n2466) );
  INVX1 U8827 ( .A(n2466), .Y(n7150) );
  AND2X1 U8828 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[28]), .Y(n2518) );
  INVX1 U8829 ( .A(n2518), .Y(n7151) );
  BUFX2 U8830 ( .A(n2305), .Y(n7152) );
  BUFX2 U8831 ( .A(n2340), .Y(n7153) );
  AND2X1 U8832 ( .A(n2271), .B(n9018), .Y(n949) );
  INVX1 U8833 ( .A(n949), .Y(n7154) );
  AND2X1 U8834 ( .A(n2247), .B(n9019), .Y(n933) );
  INVX1 U8835 ( .A(n933), .Y(n7155) );
  BUFX2 U8836 ( .A(n2380), .Y(n7156) );
  BUFX2 U8837 ( .A(n2280), .Y(n7157) );
  BUFX2 U8838 ( .A(n2356), .Y(n7158) );
  BUFX2 U8839 ( .A(n2256), .Y(n7159) );
  AND2X1 U8840 ( .A(AbeatDelay_new_reg_394[2]), .B(n9041), .Y(n2232) );
  INVX1 U8841 ( .A(n2232), .Y(n7160) );
  AND2X1 U8842 ( .A(AbeatDelay[2]), .B(n10670), .Y(n784) );
  INVX1 U8843 ( .A(n784), .Y(n7161) );
  AND2X1 U8844 ( .A(tmp_3_fu_706_p2[7]), .B(n8996), .Y(n769) );
  INVX1 U8845 ( .A(n769), .Y(n7162) );
  AND2X1 U8846 ( .A(AbeatDelay_new_reg_394[14]), .B(n9041), .Y(n2220) );
  INVX1 U8847 ( .A(n2220), .Y(n7163) );
  AND2X1 U8848 ( .A(AbeatDelay[19]), .B(n10670), .Y(n727) );
  INVX1 U8849 ( .A(n727), .Y(n7164) );
  AND2X1 U8850 ( .A(tmp_3_fu_706_p2[24]), .B(n8997), .Y(n712) );
  INVX1 U8851 ( .A(n712), .Y(n7165) );
  AND2X1 U8852 ( .A(AbeatDelay_new_reg_394[25]), .B(n9041), .Y(n2209) );
  INVX1 U8853 ( .A(n2209), .Y(n7166) );
  AND2X1 U8854 ( .A(AstimDelay[0]), .B(n10670), .Y(n684) );
  INVX1 U8855 ( .A(n684), .Y(n7167) );
  AND2X1 U8856 ( .A(tmp_6_fu_497_p3[2]), .B(n8967), .Y(n678) );
  INVX1 U8857 ( .A(n678), .Y(n7168) );
  AND2X1 U8858 ( .A(AstimDelay[17]), .B(n8896), .Y(n632) );
  INVX1 U8859 ( .A(n632), .Y(n7169) );
  AND2X1 U8860 ( .A(tmp_6_fu_497_p3[21]), .B(n8966), .Y(n621) );
  INVX1 U8861 ( .A(n621), .Y(n7170) );
  AND2X1 U8862 ( .A(VstimDelay[3]), .B(n10670), .Y(n574) );
  INVX1 U8863 ( .A(n574), .Y(n7171) );
  AND2X1 U8864 ( .A(tmp_7_fu_511_p3[9]), .B(n8965), .Y(n557) );
  INVX1 U8865 ( .A(n557), .Y(n7172) );
  AND2X1 U8866 ( .A(VstimDelay[18]), .B(n10670), .Y(n529) );
  INVX1 U8867 ( .A(n529), .Y(n7173) );
  AND2X1 U8868 ( .A(tmp_7_fu_511_p3[25]), .B(n8964), .Y(n509) );
  INVX1 U8869 ( .A(n509), .Y(n7174) );
  AND2X1 U8870 ( .A(VstimDelay[26]), .B(n10670), .Y(n505) );
  INVX1 U8871 ( .A(n505), .Y(n7175) );
  AND2X1 U8872 ( .A(\Decision_AXILiteS_s_axi_U/n360 ), .B(
        \Decision_AXILiteS_s_axi_U/n351 ), .Y(\Decision_AXILiteS_s_axi_U/n359 ) );
  INVX1 U8873 ( .A(\Decision_AXILiteS_s_axi_U/n359 ), .Y(n7176) );
  AND2X1 U8874 ( .A(\Decision_AXILiteS_s_axi_U/n356 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n409 ) );
  INVX1 U8875 ( .A(\Decision_AXILiteS_s_axi_U/n409 ), .Y(n7177) );
  AND2X1 U8876 ( .A(v_length[31]), .B(n8410), .Y(
        \Decision_AXILiteS_s_axi_U/n374 ) );
  INVX1 U8877 ( .A(\Decision_AXILiteS_s_axi_U/n374 ), .Y(n7178) );
  AND2X1 U8878 ( .A(\Decision_AXILiteS_s_axi_U/n358 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n452 ) );
  INVX1 U8879 ( .A(\Decision_AXILiteS_s_axi_U/n452 ), .Y(n7179) );
  AND2X1 U8880 ( .A(a_length[28]), .B(n8116), .Y(
        \Decision_AXILiteS_s_axi_U/n424 ) );
  INVX1 U8881 ( .A(\Decision_AXILiteS_s_axi_U/n424 ), .Y(n7180) );
  AND2X1 U8882 ( .A(\Decision_AXILiteS_s_axi_U/n364 ), .B(n8411), .Y(
        \Decision_AXILiteS_s_axi_U/n466 ) );
  INVX1 U8883 ( .A(\Decision_AXILiteS_s_axi_U/n466 ), .Y(n7181) );
  AND2X1 U8884 ( .A(vthresh[29]), .B(n7865), .Y(
        \Decision_AXILiteS_s_axi_U/n486 ) );
  INVX1 U8885 ( .A(\Decision_AXILiteS_s_axi_U/n486 ), .Y(n7182) );
  AND2X1 U8886 ( .A(s_axi_AXILiteS_AWADDR[1]), .B(n8652), .Y(
        \Decision_AXILiteS_s_axi_U/n636 ) );
  INVX1 U8887 ( .A(\Decision_AXILiteS_s_axi_U/n636 ), .Y(n7183) );
  AND2X1 U8888 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[13]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n440 )
         );
  INVX1 U8889 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n440 ), 
        .Y(n7184) );
  AND2X1 U8890 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[12]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n472 )
         );
  INVX1 U8891 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n472 ), 
        .Y(n7185) );
  AND2X1 U8892 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[15]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n512 )
         );
  INVX1 U8893 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n512 ), 
        .Y(n7186) );
  AND2X1 U8894 ( .A(n9467), .B(data_read_reg_1495[14]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n544 )
         );
  INVX1 U8895 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n544 ), 
        .Y(n7187) );
  AND2X1 U8896 ( .A(n9468), .B(data_read_reg_1495[3]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n590 )
         );
  INVX1 U8897 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n590 ), 
        .Y(n7188) );
  AND2X1 U8898 ( .A(n9468), .B(data_read_reg_1495[9]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n602 )
         );
  INVX1 U8899 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n602 ), 
        .Y(n7189) );
  AND2X1 U8900 ( .A(n9469), .B(data_read_reg_1495[2]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n622 )
         );
  INVX1 U8901 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n622 ), 
        .Y(n7190) );
  AND2X1 U8902 ( .A(n9469), .B(data_read_reg_1495[8]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n634 )
         );
  INVX1 U8903 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n634 ), 
        .Y(n7191) );
  AND2X1 U8904 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][3] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n656 )
         );
  INVX1 U8905 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n656 ), 
        .Y(n7192) );
  AND2X1 U8906 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][2] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n674 )
         );
  INVX1 U8907 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n674 ), 
        .Y(n7193) );
  AND2X1 U8908 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][1] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n691 )
         );
  INVX1 U8909 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n691 ), 
        .Y(n7194) );
  AND2X1 U8910 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][13] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n703 )
         );
  INVX1 U8911 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n703 ), 
        .Y(n7195) );
  AND2X1 U8912 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][0] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n707 )
         );
  INVX1 U8913 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n707 ), 
        .Y(n7196) );
  AND2X1 U8914 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][12] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n719 )
         );
  INVX1 U8915 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n719 ), 
        .Y(n7197) );
  AND2X1 U8916 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][15] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n739 )
         );
  INVX1 U8917 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n739 ), 
        .Y(n7198) );
  AND2X1 U8918 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][14] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n755 )
         );
  INVX1 U8919 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n755 ), 
        .Y(n7199) );
  AND2X1 U8920 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][9] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n767 )
         );
  INVX1 U8921 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n767 ), 
        .Y(n7200) );
  AND2X1 U8922 ( .A(n9466), .B(data_read_reg_1495[5]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n786 )
         );
  INVX1 U8923 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n786 ), 
        .Y(n7201) );
  AND2X1 U8924 ( .A(n9466), .B(data_read_reg_1495[11]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n798 )
         );
  INVX1 U8925 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n798 ), 
        .Y(n7202) );
  AND2X1 U8926 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][8] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n817 )
         );
  INVX1 U8927 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n817 ), 
        .Y(n7203) );
  AND2X1 U8928 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][11] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n838 )
         );
  INVX1 U8929 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n838 ), 
        .Y(n7204) );
  AND2X1 U8930 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][10] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n854 )
         );
  INVX1 U8931 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n854 ), 
        .Y(n7205) );
  AND2X1 U8932 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[4]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n870 )
         );
  INVX1 U8933 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n870 ), 
        .Y(n7206) );
  AND2X1 U8934 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[10]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n882 )
         );
  INVX1 U8935 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n882 ), 
        .Y(n7207) );
  BUFX2 U8936 ( .A(n11090), .Y(n7208) );
  AND2X1 U8937 ( .A(v_thresh[26]), .B(n9540), .Y(n12193) );
  INVX1 U8938 ( .A(n12193), .Y(n7209) );
  AND2X1 U8939 ( .A(a_thresh[26]), .B(n9490), .Y(n11560) );
  INVX1 U8940 ( .A(n11560), .Y(n7210) );
  AND2X1 U8941 ( .A(sum_reg_308[3]), .B(n8929), .Y(n2686) );
  INVX1 U8942 ( .A(n2686), .Y(n7211) );
  AND2X1 U8943 ( .A(sum_1_reg_376[1]), .B(n8930), .Y(n2412) );
  INVX1 U8944 ( .A(n2412), .Y(n7212) );
  AND2X1 U8945 ( .A(tmp_29_i_fu_752_p2[16]), .B(n8920), .Y(n3177) );
  INVX1 U8946 ( .A(n3177), .Y(n7213) );
  AND2X1 U8947 ( .A(tmp_29_i1_fu_1065_p2[16]), .B(n8922), .Y(n3229) );
  INVX1 U8948 ( .A(n3229), .Y(n7214) );
  AND2X1 U8949 ( .A(tmp_29_i_fu_752_p2[6]), .B(n8920), .Y(n3156) );
  INVX1 U8950 ( .A(n3156), .Y(n7215) );
  AND2X1 U8951 ( .A(tmp_29_i1_fu_1065_p2[6]), .B(n8922), .Y(n3208) );
  INVX1 U8952 ( .A(n3208), .Y(n7216) );
  AND2X1 U8953 ( .A(CircularBuffer_len_write_assig_fu_817_p2[10]), .B(n8894), 
        .Y(n1589) );
  INVX1 U8954 ( .A(n1589), .Y(n7217) );
  AND2X1 U8955 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[10]), .B(n8891), .Y(n913) );
  INVX1 U8956 ( .A(n913), .Y(n7218) );
  AND2X1 U8957 ( .A(sum_1_reg_376[26]), .B(n8930), .Y(n2512) );
  INVX1 U8958 ( .A(n2512), .Y(n7219) );
  AND2X1 U8959 ( .A(sum_reg_308[17]), .B(n8929), .Y(n2630) );
  INVX1 U8960 ( .A(n2630), .Y(n7220) );
  INVX1 U8961 ( .A(n4620), .Y(n7221) );
  AND2X1 U8962 ( .A(ACaptureThresh_loc_reg_288[14]), .B(n8971), .Y(n3034) );
  INVX1 U8963 ( .A(n3034), .Y(n7222) );
  BUFX2 U8964 ( .A(n3033), .Y(n7223) );
  INVX1 U8965 ( .A(n4605), .Y(n7224) );
  AND2X1 U8966 ( .A(ACaptureThresh_loc_reg_288[29]), .B(n8971), .Y(n3004) );
  INVX1 U8967 ( .A(n3004), .Y(n7225) );
  BUFX2 U8968 ( .A(n3003), .Y(n7226) );
  INVX1 U8969 ( .A(n4559), .Y(n7227) );
  AND2X1 U8970 ( .A(VCaptureThresh_loc_reg_298[11]), .B(n8970), .Y(n2912) );
  INVX1 U8971 ( .A(n2912), .Y(n7228) );
  BUFX2 U8972 ( .A(n2911), .Y(n7229) );
  INVX1 U8973 ( .A(n4544), .Y(n7230) );
  AND2X1 U8974 ( .A(VCaptureThresh_loc_reg_298[26]), .B(n8969), .Y(n2882) );
  INVX1 U8975 ( .A(n2882), .Y(n7231) );
  BUFX2 U8976 ( .A(n2881), .Y(n7232) );
  BUFX2 U8977 ( .A(n1472), .Y(n7233) );
  BUFX2 U8978 ( .A(n837), .Y(n7234) );
  AND2X1 U8979 ( .A(n1529), .B(n1530), .Y(n1520) );
  INVX1 U8980 ( .A(n1520), .Y(n7235) );
  BUFX2 U8981 ( .A(n1531), .Y(n7236) );
  AND2X1 U8982 ( .A(n807), .B(n808), .Y(n798) );
  INVX1 U8983 ( .A(n798), .Y(n7237) );
  BUFX2 U8984 ( .A(n809), .Y(n7238) );
  AND2X1 U8985 ( .A(n9921), .B(n9920), .Y(n2061) );
  INVX1 U8986 ( .A(n2061), .Y(n7239) );
  AND2X1 U8987 ( .A(recentVBools_len[2]), .B(recentVBools_len[1]), .Y(n3195)
         );
  INVX1 U8988 ( .A(n3195), .Y(n7240) );
  AND2X1 U8989 ( .A(recentABools_len[2]), .B(recentABools_len[1]), .Y(n3247)
         );
  INVX1 U8990 ( .A(n3247), .Y(n7241) );
  AND2X1 U8991 ( .A(n10506), .B(n10510), .Y(n319) );
  INVX1 U8992 ( .A(n319), .Y(n7242) );
  AND2X1 U8993 ( .A(n9866), .B(n9865), .Y(n1951) );
  INVX1 U8994 ( .A(n1951), .Y(n7243) );
  AND2X1 U8995 ( .A(n10713), .B(n10715), .Y(n282) );
  INVX1 U8996 ( .A(n282), .Y(n7244) );
  AND2X1 U8997 ( .A(n9851), .B(n9852), .Y(n2047) );
  INVX1 U8998 ( .A(n2047), .Y(n7245) );
  AND2X1 U8999 ( .A(n8660), .B(n9961), .Y(n1817) );
  INVX1 U9000 ( .A(n1817), .Y(n7246) );
  AND2X1 U9001 ( .A(n9937), .B(n9936), .Y(n1818) );
  INVX1 U9002 ( .A(n1818), .Y(n7247) );
  BUFX2 U9003 ( .A(n1816), .Y(n7248) );
  AND2X1 U9004 ( .A(n8661), .B(n10269), .Y(n1255) );
  INVX1 U9005 ( .A(n1255), .Y(n7249) );
  AND2X1 U9006 ( .A(n10245), .B(n10244), .Y(n1256) );
  INVX1 U9007 ( .A(n1256), .Y(n7250) );
  BUFX2 U9008 ( .A(n1254), .Y(n7251) );
  INVX1 U9009 ( .A(recentABools_data_address0[0]), .Y(n7252) );
  BUFX2 U9010 ( .A(n395), .Y(n7253) );
  BUFX2 U9011 ( .A(n394), .Y(n7254) );
  AND2X1 U9012 ( .A(recentdatapoints_len_load_op_fu_556_p2[8]), .B(n8972), .Y(
        n1828) );
  INVX1 U9013 ( .A(n1828), .Y(n7255) );
  AND2X1 U9014 ( .A(recentdatapoints_len_load_op_fu_556_p2[22]), .B(n8972), 
        .Y(n1847) );
  INVX1 U9015 ( .A(n1847), .Y(n7256) );
  AND2X1 U9016 ( .A(p_tmp_i_fu_587_p3[3]), .B(n8975), .Y(n1867) );
  INVX1 U9017 ( .A(n1867), .Y(n7257) );
  AND2X1 U9018 ( .A(n10895), .B(n10897), .Y(\Decision_AXILiteS_s_axi_U/n481 )
         );
  INVX1 U9019 ( .A(\Decision_AXILiteS_s_axi_U/n481 ), .Y(n7258) );
  AND2X1 U9020 ( .A(CircularBuffer_len_read_assign_fu_772_p2[30]), .B(n3151), 
        .Y(n2734) );
  INVX1 U9021 ( .A(n2734), .Y(n7259) );
  AND2X1 U9022 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[30]), .B(n3149), .Y(n2238) );
  INVX1 U9023 ( .A(n2238), .Y(n7260) );
  AND2X1 U9024 ( .A(recentdatapoints_data_q0[2]), .B(n8869), .Y(n414) );
  INVX1 U9025 ( .A(n414), .Y(n7261) );
  AND2X1 U9026 ( .A(recentdatapoints_data_q0[11]), .B(n8868), .Y(n425) );
  INVX1 U9027 ( .A(n425), .Y(n7262) );
  AND2X1 U9028 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[9]), 
        .Y(n442) );
  INVX1 U9029 ( .A(n442), .Y(n7263) );
  AND2X1 U9030 ( .A(CircularBuffer_len_read_assign_fu_772_p2[21]), .B(n8919), 
        .Y(n2752) );
  INVX1 U9031 ( .A(n2752), .Y(n7264) );
  AND2X1 U9032 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[21]), .B(n8921), .Y(n2259) );
  INVX1 U9033 ( .A(n2259), .Y(n7265) );
  AND2X1 U9034 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n71 ), .B(n8887), .Y(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n48 ) );
  INVX1 U9035 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n48 ), 
        .Y(n7266) );
  AND2X1 U9036 ( .A(n4694), .B(\tmp_12_reg_1694[0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n77 ) );
  INVX1 U9037 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n77 ), 
        .Y(n7267) );
  AND2X1 U9038 ( .A(n8882), .B(\Decision_AXILiteS_s_axi_U/n396 ), .Y(
        \Decision_AXILiteS_s_axi_U/n495 ) );
  INVX1 U9039 ( .A(\Decision_AXILiteS_s_axi_U/n495 ), .Y(n7268) );
  AND2X1 U9040 ( .A(\Decision_AXILiteS_s_axi_U/n533 ), .B(
        \Decision_AXILiteS_s_axi_U/n352 ), .Y(\Decision_AXILiteS_s_axi_U/n547 ) );
  INVX1 U9041 ( .A(\Decision_AXILiteS_s_axi_U/n547 ), .Y(n7269) );
  BUFX2 U9042 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n32 ), 
        .Y(n7270) );
  AND2X1 U9043 ( .A(a_length[10]), .B(n8952), .Y(n3106) );
  INVX1 U9044 ( .A(n3106), .Y(n7271) );
  AND2X1 U9045 ( .A(a_length[28]), .B(n8953), .Y(n3070) );
  INVX1 U9046 ( .A(n3070), .Y(n7272) );
  AND2X1 U9047 ( .A(v_length[20]), .B(n8955), .Y(n2958) );
  INVX1 U9048 ( .A(n2958), .Y(n7273) );
  AND2X1 U9049 ( .A(v_length[30]), .B(n8954), .Y(n2938) );
  INVX1 U9050 ( .A(n2938), .Y(n7274) );
  AND2X1 U9051 ( .A(recentdatapoints_head_i[16]), .B(n8980), .Y(n1967) );
  INVX1 U9052 ( .A(n1967), .Y(n7275) );
  AND2X1 U9053 ( .A(recentdatapoints_head_i[27]), .B(n8979), .Y(n1956) );
  INVX1 U9054 ( .A(n1956), .Y(n7276) );
  AND2X1 U9055 ( .A(p_tmp_i_reg_1556[20]), .B(n8979), .Y(n1902) );
  INVX1 U9056 ( .A(n1902), .Y(n7277) );
  AND2X1 U9057 ( .A(p_tmp_i_reg_1556[9]), .B(n8978), .Y(n1880) );
  INVX1 U9058 ( .A(n1880), .Y(n7278) );
  AND2X1 U9059 ( .A(ap_CS_fsm[2]), .B(recentVBools_head_i[3]), .Y(n1798) );
  INVX1 U9060 ( .A(n1798), .Y(n7279) );
  AND2X1 U9061 ( .A(recentVBools_head_i[24]), .B(n9009), .Y(n1732) );
  INVX1 U9062 ( .A(n1732), .Y(n7280) );
  AND2X1 U9063 ( .A(n2768), .B(n8992), .Y(n1629) );
  INVX1 U9064 ( .A(n1629), .Y(n7281) );
  AND2X1 U9065 ( .A(n2748), .B(n8991), .Y(n1616) );
  INVX1 U9066 ( .A(n1616), .Y(n7282) );
  BUFX2 U9067 ( .A(n2781), .Y(n7283) );
  BUFX2 U9068 ( .A(n2765), .Y(n7284) );
  BUFX2 U9069 ( .A(n2817), .Y(n7285) );
  AND2X1 U9070 ( .A(CircularBuffer_len_write_assig_fu_817_p2[9]), .B(n8894), 
        .Y(n1590) );
  INVX1 U9071 ( .A(n1590), .Y(n7286) );
  AND2X1 U9072 ( .A(CircularBuffer_sum_read_assign_reg_1610[18]), .B(n9005), 
        .Y(n1430) );
  INVX1 U9073 ( .A(n1430), .Y(n7287) );
  AND2X1 U9074 ( .A(CircularBuffer_sum_read_assign_reg_1610[22]), .B(n9007), 
        .Y(n1422) );
  INVX1 U9075 ( .A(n1422), .Y(n7288) );
  AND2X1 U9076 ( .A(CircularBuffer_sum_read_assign_reg_1610[24]), .B(n9006), 
        .Y(n1418) );
  INVX1 U9077 ( .A(n1418), .Y(n7289) );
  BUFX2 U9078 ( .A(n2731), .Y(n7290) );
  BUFX2 U9079 ( .A(n2719), .Y(n7291) );
  AND2X1 U9080 ( .A(n9012), .B(sum_phi_fu_311_p4[14]), .Y(n2640) );
  INVX1 U9081 ( .A(n2640), .Y(n7292) );
  BUFX2 U9082 ( .A(n2705), .Y(n7293) );
  AND2X1 U9083 ( .A(n9012), .B(sum_phi_fu_311_p4[30]), .Y(n2576) );
  INVX1 U9084 ( .A(n2576), .Y(n7294) );
  AND2X1 U9085 ( .A(recentABools_head_i[11]), .B(n9040), .Y(n1316) );
  INVX1 U9086 ( .A(n1316), .Y(n7295) );
  AND2X1 U9087 ( .A(recentABools_head_i[22]), .B(n9039), .Y(n1291) );
  INVX1 U9088 ( .A(n1291), .Y(n7296) );
  AND2X1 U9089 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[28]), .B(n9038), 
        .Y(n1277) );
  INVX1 U9090 ( .A(n1277), .Y(n7297) );
  AND2X1 U9091 ( .A(recentABools_head_i[4]), .B(ap_CS_fsm[7]), .Y(n1226) );
  INVX1 U9092 ( .A(n1226), .Y(n7298) );
  AND2X1 U9093 ( .A(VbeatFallDelay[10]), .B(n9036), .Y(n1166) );
  INVX1 U9094 ( .A(n1166), .Y(n7299) );
  AND2X1 U9095 ( .A(VbeatFallDelay_new_1_reg_342[13]), .B(n9013), .Y(n2170) );
  INVX1 U9096 ( .A(n2170), .Y(n7300) );
  AND2X1 U9097 ( .A(tmp_5_fu_726_p2[14]), .B(n8993), .Y(n1152) );
  INVX1 U9098 ( .A(n1152), .Y(n7301) );
  AND2X1 U9099 ( .A(VbeatFallDelay[21]), .B(n9035), .Y(n1122) );
  INVX1 U9100 ( .A(n1122), .Y(n7302) );
  AND2X1 U9101 ( .A(VbeatFallDelay_new_1_reg_342[27]), .B(n9013), .Y(n2184) );
  INVX1 U9102 ( .A(n2184), .Y(n7303) );
  AND2X1 U9103 ( .A(VbeatFallDelay[31]), .B(n9034), .Y(n1082) );
  INVX1 U9104 ( .A(n1082), .Y(n7304) );
  AND2X1 U9105 ( .A(n10452), .B(n8994), .Y(n1078) );
  INVX1 U9106 ( .A(n1078), .Y(n7305) );
  AND2X1 U9107 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[4]), .Y(n2562) );
  INVX1 U9108 ( .A(n2562), .Y(n7306) );
  AND2X1 U9109 ( .A(VbeatDelay[12]), .B(n9032), .Y(n1037) );
  INVX1 U9110 ( .A(n1037), .Y(n7307) );
  AND2X1 U9111 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[17]), .Y(n2549) );
  INVX1 U9112 ( .A(n2549), .Y(n7308) );
  AND2X1 U9113 ( .A(tmp_4_fu_716_p2[19]), .B(n8995), .Y(n1016) );
  INVX1 U9114 ( .A(n1016), .Y(n7309) );
  AND2X1 U9115 ( .A(VbeatDelay[21]), .B(n9031), .Y(n1007) );
  INVX1 U9116 ( .A(n1007), .Y(n7310) );
  AND2X1 U9117 ( .A(VbeatDelay[26]), .B(n9033), .Y(n990) );
  INVX1 U9118 ( .A(n990), .Y(n7311) );
  AND2X1 U9119 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[28]), .Y(n2538) );
  INVX1 U9120 ( .A(n2538), .Y(n7312) );
  BUFX2 U9121 ( .A(n2323), .Y(n7313) );
  AND2X1 U9122 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[17]), .Y(n2474) );
  INVX1 U9123 ( .A(n2474), .Y(n7314) );
  BUFX2 U9124 ( .A(n2310), .Y(n7315) );
  AND2X1 U9125 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[29]), .Y(n2522) );
  INVX1 U9126 ( .A(n2522), .Y(n7316) );
  AND2X1 U9127 ( .A(n2281), .B(n9019), .Y(n957) );
  INVX1 U9128 ( .A(n957), .Y(n7317) );
  AND2X1 U9129 ( .A(n2255), .B(n9018), .Y(n940) );
  INVX1 U9130 ( .A(n940), .Y(n7318) );
  BUFX2 U9131 ( .A(n2294), .Y(n7319) );
  BUFX2 U9132 ( .A(n2382), .Y(n7320) );
  BUFX2 U9133 ( .A(n2272), .Y(n7321) );
  BUFX2 U9134 ( .A(n2354), .Y(n7322) );
  BUFX2 U9135 ( .A(n2248), .Y(n7323) );
  BUFX2 U9136 ( .A(n2344), .Y(n7324) );
  AND2X1 U9137 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[9]), .B(n8891), 
        .Y(n914) );
  INVX1 U9138 ( .A(n914), .Y(n7325) );
  AND2X1 U9139 ( .A(AbeatDelay_new_reg_394[3]), .B(n9041), .Y(n2231) );
  INVX1 U9140 ( .A(n2231), .Y(n7326) );
  AND2X1 U9141 ( .A(tmp_3_fu_706_p2[8]), .B(n8996), .Y(n766) );
  INVX1 U9142 ( .A(n766), .Y(n7327) );
  AND2X1 U9143 ( .A(AbeatDelay_new_reg_394[15]), .B(n9041), .Y(n2219) );
  INVX1 U9144 ( .A(n2219), .Y(n7328) );
  AND2X1 U9145 ( .A(AbeatDelay[20]), .B(n10670), .Y(n723) );
  INVX1 U9146 ( .A(n723), .Y(n7329) );
  AND2X1 U9147 ( .A(AbeatDelay_new_reg_394[26]), .B(n9041), .Y(n2208) );
  INVX1 U9148 ( .A(n2208), .Y(n7330) );
  AND2X1 U9149 ( .A(tmp_3_fu_706_p2[27]), .B(n8997), .Y(n702) );
  INVX1 U9150 ( .A(n702), .Y(n7331) );
  AND2X1 U9151 ( .A(AstimDelay[1]), .B(n10670), .Y(n680) );
  INVX1 U9152 ( .A(n680), .Y(n7332) );
  AND2X1 U9153 ( .A(AstimDelay[18]), .B(n8896), .Y(n629) );
  INVX1 U9154 ( .A(n629), .Y(n7333) );
  AND2X1 U9155 ( .A(tmp_6_fu_497_p3[22]), .B(n8966), .Y(n618) );
  INVX1 U9156 ( .A(n618), .Y(n7334) );
  AND2X1 U9157 ( .A(VstimDelay[4]), .B(n8896), .Y(n571) );
  INVX1 U9158 ( .A(n571), .Y(n7335) );
  AND2X1 U9159 ( .A(tmp_7_fu_511_p3[7]), .B(n8965), .Y(n563) );
  INVX1 U9160 ( .A(n563), .Y(n7336) );
  AND2X1 U9161 ( .A(VstimDelay[19]), .B(n10670), .Y(n526) );
  INVX1 U9162 ( .A(n526), .Y(n7337) );
  AND2X1 U9163 ( .A(tmp_7_fu_511_p3[23]), .B(n8963), .Y(n515) );
  INVX1 U9164 ( .A(n515), .Y(n7338) );
  AND2X1 U9165 ( .A(tmp_7_fu_511_p3[26]), .B(n8964), .Y(n506) );
  INVX1 U9166 ( .A(n506), .Y(n7339) );
  AND2X1 U9167 ( .A(VstimDelay[27]), .B(n10670), .Y(n502) );
  INVX1 U9168 ( .A(n502), .Y(n7340) );
  AND2X1 U9169 ( .A(v_length[29]), .B(n8410), .Y(
        \Decision_AXILiteS_s_axi_U/n377 ) );
  INVX1 U9170 ( .A(\Decision_AXILiteS_s_axi_U/n377 ), .Y(n7341) );
  AND2X1 U9171 ( .A(\Decision_AXILiteS_s_axi_U/n356 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n451 ) );
  INVX1 U9172 ( .A(\Decision_AXILiteS_s_axi_U/n451 ), .Y(n7342) );
  AND2X1 U9173 ( .A(a_length[31]), .B(n8116), .Y(
        \Decision_AXILiteS_s_axi_U/n420 ) );
  INVX1 U9174 ( .A(\Decision_AXILiteS_s_axi_U/n420 ), .Y(n7343) );
  AND2X1 U9175 ( .A(\Decision_AXILiteS_s_axi_U/n362 ), .B(n8411), .Y(
        \Decision_AXILiteS_s_axi_U/n465 ) );
  INVX1 U9176 ( .A(\Decision_AXILiteS_s_axi_U/n465 ), .Y(n7344) );
  AND2X1 U9177 ( .A(vthresh[30]), .B(n7865), .Y(
        \Decision_AXILiteS_s_axi_U/n485 ) );
  INVX1 U9178 ( .A(\Decision_AXILiteS_s_axi_U/n485 ), .Y(n7345) );
  AND2X1 U9179 ( .A(s_axi_AXILiteS_AWADDR[2]), .B(n8652), .Y(
        \Decision_AXILiteS_s_axi_U/n637 ) );
  INVX1 U9180 ( .A(\Decision_AXILiteS_s_axi_U/n637 ), .Y(n7346) );
  AND2X1 U9181 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[12]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n438 )
         );
  INVX1 U9182 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n438 ), 
        .Y(n7347) );
  AND2X1 U9183 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[13]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n474 )
         );
  INVX1 U9184 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n474 ), 
        .Y(n7348) );
  AND2X1 U9185 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[14]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n510 )
         );
  INVX1 U9186 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n510 ), 
        .Y(n7349) );
  AND2X1 U9187 ( .A(n9467), .B(data_read_reg_1495[15]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n546 )
         );
  INVX1 U9188 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n546 ), 
        .Y(n7350) );
  AND2X1 U9189 ( .A(n9468), .B(data_read_reg_1495[2]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n588 )
         );
  INVX1 U9190 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n588 ), 
        .Y(n7351) );
  AND2X1 U9191 ( .A(n9468), .B(data_read_reg_1495[8]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n600 )
         );
  INVX1 U9192 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n600 ), 
        .Y(n7352) );
  AND2X1 U9193 ( .A(n9469), .B(data_read_reg_1495[3]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n624 )
         );
  INVX1 U9194 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n624 ), 
        .Y(n7353) );
  AND2X1 U9195 ( .A(n9469), .B(data_read_reg_1495[9]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n636 )
         );
  INVX1 U9196 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n636 ), 
        .Y(n7354) );
  AND2X1 U9197 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][2] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n655 )
         );
  INVX1 U9198 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n655 ), 
        .Y(n7355) );
  AND2X1 U9199 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][3] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n675 )
         );
  INVX1 U9200 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n675 ), 
        .Y(n7356) );
  AND2X1 U9201 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][0] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n690 )
         );
  INVX1 U9202 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n690 ), 
        .Y(n7357) );
  AND2X1 U9203 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][12] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n702 )
         );
  INVX1 U9204 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n702 ), 
        .Y(n7358) );
  AND2X1 U9205 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][1] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n708 )
         );
  INVX1 U9206 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n708 ), 
        .Y(n7359) );
  AND2X1 U9207 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][13] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n720 )
         );
  INVX1 U9208 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n720 ), 
        .Y(n7360) );
  AND2X1 U9209 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][14] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n738 )
         );
  INVX1 U9210 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n738 ), 
        .Y(n7361) );
  AND2X1 U9211 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][15] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n756 )
         );
  INVX1 U9212 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n756 ), 
        .Y(n7362) );
  AND2X1 U9213 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][8] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n766 )
         );
  INVX1 U9214 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n766 ), 
        .Y(n7363) );
  AND2X1 U9215 ( .A(n9466), .B(data_read_reg_1495[4]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n784 )
         );
  INVX1 U9216 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n784 ), 
        .Y(n7364) );
  AND2X1 U9217 ( .A(n9466), .B(data_read_reg_1495[10]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n796 )
         );
  INVX1 U9218 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n796 ), 
        .Y(n7365) );
  AND2X1 U9219 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][9] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n818 )
         );
  INVX1 U9220 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n818 ), 
        .Y(n7366) );
  AND2X1 U9221 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][10] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n837 )
         );
  INVX1 U9222 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n837 ), 
        .Y(n7367) );
  AND2X1 U9223 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][11] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n855 )
         );
  INVX1 U9224 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n855 ), 
        .Y(n7368) );
  AND2X1 U9225 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[5]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n872 )
         );
  INVX1 U9226 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n872 ), 
        .Y(n7369) );
  AND2X1 U9227 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[11]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n884 )
         );
  INVX1 U9228 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n884 ), 
        .Y(n7370) );
  AND2X1 U9229 ( .A(tmp_29_i_fu_752_p2[15]), .B(n8920), .Y(n3178) );
  INVX1 U9230 ( .A(n3178), .Y(n7371) );
  AND2X1 U9231 ( .A(tmp_29_i1_fu_1065_p2[15]), .B(n8922), .Y(n3230) );
  INVX1 U9232 ( .A(n3230), .Y(n7372) );
  AND2X1 U9233 ( .A(tmp_29_i_fu_752_p2[5]), .B(n8920), .Y(n3157) );
  INVX1 U9234 ( .A(n3157), .Y(n7373) );
  AND2X1 U9235 ( .A(tmp_29_i1_fu_1065_p2[5]), .B(n8922), .Y(n3209) );
  INVX1 U9236 ( .A(n3209), .Y(n7374) );
  AND2X1 U9237 ( .A(ap_rst_n), .B(\Decision_AXILiteS_s_axi_U/n602 ), .Y(
        \Decision_AXILiteS_s_axi_U/n601 ) );
  INVX1 U9238 ( .A(\Decision_AXILiteS_s_axi_U/n601 ), .Y(n7375) );
  AND2X1 U9239 ( .A(sum_reg_308[21]), .B(n8929), .Y(n2614) );
  INVX1 U9240 ( .A(n2614), .Y(n7376) );
  AND2X1 U9241 ( .A(sum_1_reg_376[25]), .B(n8930), .Y(n2508) );
  INVX1 U9242 ( .A(n2508), .Y(n7377) );
  AND2X1 U9243 ( .A(sum_1_reg_376[2]), .B(n8930), .Y(n2416) );
  INVX1 U9244 ( .A(n2416), .Y(n7378) );
  AND2X1 U9245 ( .A(sum_reg_308[16]), .B(n8929), .Y(n2634) );
  INVX1 U9246 ( .A(n2634), .Y(n7379) );
  AND2X1 U9247 ( .A(datapointV_1_fu_674_p2[16]), .B(n397), .Y(n399) );
  INVX1 U9248 ( .A(n399), .Y(n7380) );
  AND2X1 U9249 ( .A(datapointA_1_fu_1017_p2[16]), .B(n439), .Y(n441) );
  INVX1 U9250 ( .A(n441), .Y(n7381) );
  INVX1 U9251 ( .A(n3858), .Y(n7382) );
  AND2X1 U9252 ( .A(CircularBuffer_head_i_read_ass_reg_1624[3]), .B(n9008), 
        .Y(n1704) );
  INVX1 U9253 ( .A(n1704), .Y(n7383) );
  INVX1 U9254 ( .A(n3659), .Y(n7384) );
  AND2X1 U9255 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[4]), .B(n9037), 
        .Y(n1229) );
  INVX1 U9256 ( .A(n1229), .Y(n7385) );
  INVX1 U9257 ( .A(n4619), .Y(n7386) );
  AND2X1 U9258 ( .A(ACaptureThresh_loc_reg_288[15]), .B(n8968), .Y(n3032) );
  INVX1 U9259 ( .A(n3032), .Y(n7387) );
  BUFX2 U9260 ( .A(n3031), .Y(n7388) );
  INVX1 U9261 ( .A(n4604), .Y(n7389) );
  AND2X1 U9262 ( .A(ACaptureThresh_loc_reg_288[30]), .B(n8971), .Y(n3002) );
  INVX1 U9263 ( .A(n3002), .Y(n7390) );
  BUFX2 U9264 ( .A(n3001), .Y(n7391) );
  INVX1 U9265 ( .A(n4558), .Y(n7392) );
  AND2X1 U9266 ( .A(VCaptureThresh_loc_reg_298[12]), .B(n8970), .Y(n2910) );
  INVX1 U9267 ( .A(n2910), .Y(n7393) );
  BUFX2 U9268 ( .A(n2909), .Y(n7394) );
  INVX1 U9269 ( .A(n4543), .Y(n7395) );
  AND2X1 U9270 ( .A(VCaptureThresh_loc_reg_298[27]), .B(n8969), .Y(n2880) );
  INVX1 U9271 ( .A(n2880), .Y(n7396) );
  BUFX2 U9272 ( .A(n2879), .Y(n7397) );
  AND2X1 U9273 ( .A(\recentABools_data_q1[0] ), .B(n10534), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n3 ) );
  INVX1 U9274 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n3 ), 
        .Y(n7398) );
  BUFX2 U9275 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n1 ), 
        .Y(n7399) );
  BUFX2 U9276 ( .A(n12103), .Y(n7400) );
  AND2X1 U9277 ( .A(n2776), .B(n9677), .Y(n12102) );
  INVX1 U9278 ( .A(n12102), .Y(n7401) );
  BUFX2 U9279 ( .A(n11639), .Y(n7402) );
  AND2X1 U9280 ( .A(n2283), .B(n9573), .Y(n11638) );
  INVX1 U9281 ( .A(n11638), .Y(n7403) );
  BUFX2 U9282 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n26 ), 
        .Y(n7404) );
  OR2X1 U9283 ( .A(recentVBools_data_address0[1]), .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n117 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n121 ) );
  INVX1 U9284 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n121 ), .Y(n7405) );
  BUFX2 U9285 ( .A(n11166), .Y(n7406) );
  BUFX2 U9286 ( .A(n11164), .Y(n7407) );
  AND2X1 U9287 ( .A(n9905), .B(n9904), .Y(n1686) );
  INVX1 U9288 ( .A(n1686), .Y(n7408) );
  AND2X1 U9289 ( .A(n10089), .B(n10090), .Y(n1489) );
  INVX1 U9290 ( .A(n1489), .Y(n7409) );
  AND2X1 U9291 ( .A(n10584), .B(n10585), .Y(n854) );
  INVX1 U9292 ( .A(n854), .Y(n7410) );
  AND2X1 U9293 ( .A(n1547), .B(n1548), .Y(n1538) );
  INVX1 U9294 ( .A(n1538), .Y(n7411) );
  AND2X1 U9295 ( .A(n10153), .B(n10154), .Y(n1549) );
  INVX1 U9296 ( .A(n1549), .Y(n7412) );
  AND2X1 U9297 ( .A(n825), .B(n826), .Y(n816) );
  INVX1 U9298 ( .A(n816), .Y(n7413) );
  AND2X1 U9299 ( .A(n10648), .B(n10649), .Y(n827) );
  INVX1 U9300 ( .A(n827), .Y(n7414) );
  AND2X1 U9301 ( .A(n10677), .B(n10699), .Y(n272) );
  INVX1 U9302 ( .A(n272), .Y(n7415) );
  AND2X1 U9303 ( .A(n10120), .B(n10121), .Y(n3194) );
  INVX1 U9304 ( .A(n3194), .Y(n7416) );
  AND2X1 U9305 ( .A(n10615), .B(n10616), .Y(n3246) );
  INVX1 U9306 ( .A(n3246), .Y(n7417) );
  AND2X1 U9307 ( .A(n9917), .B(n9916), .Y(n2060) );
  INVX1 U9308 ( .A(n2060), .Y(n7418) );
  AND2X1 U9309 ( .A(n9831), .B(n9833), .Y(n2043) );
  INVX1 U9310 ( .A(n2043), .Y(n7419) );
  AND2X1 U9311 ( .A(n9857), .B(n9858), .Y(n2044) );
  INVX1 U9312 ( .A(n2044), .Y(n7420) );
  BUFX2 U9313 ( .A(n2042), .Y(n7421) );
  AND2X1 U9314 ( .A(n9951), .B(n9950), .Y(n1807) );
  INVX1 U9315 ( .A(n1807), .Y(n7422) );
  AND2X1 U9316 ( .A(n9953), .B(n9952), .Y(n1808) );
  INVX1 U9317 ( .A(n1808), .Y(n7423) );
  BUFX2 U9318 ( .A(n1806), .Y(n7424) );
  AND2X1 U9319 ( .A(n10259), .B(n10258), .Y(n1237) );
  INVX1 U9320 ( .A(n1237), .Y(n7425) );
  AND2X1 U9321 ( .A(n10261), .B(n10260), .Y(n1238) );
  INVX1 U9322 ( .A(n1238), .Y(n7426) );
  BUFX2 U9323 ( .A(n1236), .Y(n7427) );
  INVX1 U9324 ( .A(recentVBools_data_address0[0]), .Y(n7428) );
  BUFX2 U9325 ( .A(n381), .Y(n7429) );
  BUFX2 U9326 ( .A(n380), .Y(n7430) );
  AND2X1 U9327 ( .A(recentdatapoints_len_load_op_fu_556_p2[9]), .B(n8972), .Y(
        n1829) );
  INVX1 U9328 ( .A(n1829), .Y(n7431) );
  AND2X1 U9329 ( .A(recentdatapoints_len_load_op_fu_556_p2[23]), .B(n8972), 
        .Y(n1848) );
  INVX1 U9330 ( .A(n1848), .Y(n7432) );
  BUFX2 U9331 ( .A(n1869), .Y(n7433) );
  BUFX2 U9332 ( .A(\Decision_AXILiteS_s_axi_U/n418 ), .Y(n7434) );
  AND2X1 U9333 ( .A(n8382), .B(ap_rst_n), .Y(\Decision_AXILiteS_s_axi_U/n371 )
         );
  AND2X1 U9334 ( .A(recentdatapoints_data_q0[6]), .B(n8869), .Y(n406) );
  INVX1 U9335 ( .A(n406), .Y(n7435) );
  AND2X1 U9336 ( .A(recentdatapoints_data_q0[8]), .B(n8868), .Y(n402) );
  INVX1 U9337 ( .A(n402), .Y(n7436) );
  AND2X1 U9338 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[5]), 
        .Y(n450) );
  INVX1 U9339 ( .A(n450), .Y(n7437) );
  AND2X1 U9340 ( .A(CircularBuffer_len_read_assign_fu_772_p2[12]), .B(n3151), 
        .Y(n2770) );
  INVX1 U9341 ( .A(n2770), .Y(n7438) );
  AND2X1 U9342 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[12]), .B(n3149), .Y(n2277) );
  INVX1 U9343 ( .A(n2277), .Y(n7439) );
  AND2X1 U9344 ( .A(CircularBuffer_len_read_assign_fu_772_p2[5]), .B(n3151), 
        .Y(n2784) );
  INVX1 U9345 ( .A(n2784), .Y(n7440) );
  AND2X1 U9346 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[5]), .B(n3149), 
        .Y(n2291) );
  INVX1 U9347 ( .A(n2291), .Y(n7441) );
  AND2X1 U9348 ( .A(CircularBuffer_len_read_assign_fu_772_p2[18]), .B(n8919), 
        .Y(n2758) );
  INVX1 U9349 ( .A(n2758), .Y(n7442) );
  AND2X1 U9350 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[18]), .B(n8921), .Y(n2265) );
  INVX1 U9351 ( .A(n2265), .Y(n7443) );
  AND2X1 U9352 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n73 ), .B(n8885), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n50 ) );
  INVX1 U9353 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n50 ), 
        .Y(n7444) );
  AND2X1 U9354 ( .A(recentABools_data_address0[1]), .B(n7648), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n73 ) );
  AND2X1 U9355 ( .A(n8882), .B(\Decision_AXILiteS_s_axi_U/n352 ), .Y(
        \Decision_AXILiteS_s_axi_U/n505 ) );
  INVX1 U9356 ( .A(\Decision_AXILiteS_s_axi_U/n505 ), .Y(n7445) );
  AND2X1 U9357 ( .A(\Decision_AXILiteS_s_axi_U/n533 ), .B(
        \Decision_AXILiteS_s_axi_U/n396 ), .Y(\Decision_AXILiteS_s_axi_U/n537 ) );
  INVX1 U9358 ( .A(\Decision_AXILiteS_s_axi_U/n537 ), .Y(n7446) );
  AND2X1 U9359 ( .A(\Decision_AXILiteS_s_axi_U/n353 ), .B(
        \Decision_AXILiteS_s_axi_U/n351 ), .Y(\Decision_AXILiteS_s_axi_U/n341 ) );
  INVX1 U9360 ( .A(\Decision_AXILiteS_s_axi_U/n341 ), .Y(n7447) );
  BUFX2 U9361 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n34 ), 
        .Y(n7448) );
  AND2X1 U9362 ( .A(n9932), .B(\tmp_s_reg_1578[0] ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n33 ) );
  INVX1 U9363 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n33 ), 
        .Y(n7449) );
  OR2X1 U9364 ( .A(CircularBuffer_len_read_assign_3_reg_1711[30]), .B(n8833), 
        .Y(n8852) );
  OR2X1 U9365 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[30] ), .B(n8633), .Y(n8847) );
  AND2X1 U9366 ( .A(v_flip[0]), .B(n8951), .Y(n3138) );
  INVX1 U9367 ( .A(n3138), .Y(n7450) );
  AND2X1 U9368 ( .A(a_length[11]), .B(n8952), .Y(n3104) );
  INVX1 U9369 ( .A(n3104), .Y(n7451) );
  AND2X1 U9370 ( .A(a_length[29]), .B(n8953), .Y(n3068) );
  INVX1 U9371 ( .A(n3068), .Y(n7452) );
  AND2X1 U9372 ( .A(v_length[21]), .B(n8955), .Y(n2956) );
  INVX1 U9373 ( .A(n2956), .Y(n7453) );
  AND2X1 U9374 ( .A(v_length[31]), .B(n8954), .Y(n2936) );
  INVX1 U9375 ( .A(n2936), .Y(n7454) );
  AND2X1 U9376 ( .A(recentdatapoints_head_i[17]), .B(n8980), .Y(n1966) );
  INVX1 U9377 ( .A(n1966), .Y(n7455) );
  AND2X1 U9378 ( .A(recentdatapoints_head_i[28]), .B(n8979), .Y(n1955) );
  INVX1 U9379 ( .A(n1955), .Y(n7456) );
  AND2X1 U9380 ( .A(p_tmp_i_reg_1556[22]), .B(n8979), .Y(n1906) );
  INVX1 U9381 ( .A(n1906), .Y(n7457) );
  AND2X1 U9382 ( .A(p_tmp_i_reg_1556[8]), .B(n8979), .Y(n1878) );
  INVX1 U9383 ( .A(n1878), .Y(n7458) );
  AND2X1 U9384 ( .A(ap_CS_fsm[2]), .B(recentVBools_head_i[0]), .Y(n1792) );
  INVX1 U9385 ( .A(n1792), .Y(n7459) );
  AND2X1 U9386 ( .A(CircularBuffer_head_i_read_ass_reg_1624[25]), .B(n9009), 
        .Y(n1730) );
  INVX1 U9387 ( .A(n1730), .Y(n7460) );
  AND2X1 U9388 ( .A(n2862), .B(n8991), .Y(n1603) );
  INVX1 U9389 ( .A(n1603), .Y(n7461) );
  BUFX2 U9390 ( .A(n2779), .Y(n7462) );
  BUFX2 U9391 ( .A(n2757), .Y(n7463) );
  BUFX2 U9392 ( .A(n2821), .Y(n7464) );
  AND2X1 U9393 ( .A(CircularBuffer_len_write_assig_fu_817_p2[23]), .B(n1646), 
        .Y(n1568) );
  INVX1 U9394 ( .A(n1568), .Y(n7465) );
  AND2X1 U9395 ( .A(CircularBuffer_sum_read_assign_reg_1610[19]), .B(n9005), 
        .Y(n1428) );
  INVX1 U9396 ( .A(n1428), .Y(n7466) );
  AND2X1 U9397 ( .A(CircularBuffer_sum_read_assign_reg_1610[23]), .B(n9006), 
        .Y(n1420) );
  INVX1 U9398 ( .A(n1420), .Y(n7467) );
  AND2X1 U9399 ( .A(CircularBuffer_sum_read_assign_reg_1610[27]), .B(n9007), 
        .Y(n1412) );
  INVX1 U9400 ( .A(n1412), .Y(n7468) );
  BUFX2 U9401 ( .A(n2730), .Y(n7469) );
  AND2X1 U9402 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[13]), .Y(n2644) );
  INVX1 U9403 ( .A(n2644), .Y(n7470) );
  BUFX2 U9404 ( .A(n2717), .Y(n7471) );
  AND2X1 U9405 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[28]), .Y(n2584) );
  INVX1 U9406 ( .A(n2584), .Y(n7472) );
  BUFX2 U9407 ( .A(n2704), .Y(n7473) );
  AND2X1 U9408 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[24]), .B(n9031), 
        .Y(n1388) );
  INVX1 U9409 ( .A(n1388), .Y(n7474) );
  AND2X1 U9410 ( .A(recentABools_head_i[17]), .B(n9040), .Y(n1304) );
  INVX1 U9411 ( .A(n1304), .Y(n7475) );
  AND2X1 U9412 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[23]), .B(n9039), 
        .Y(n1289) );
  INVX1 U9413 ( .A(n1289), .Y(n7476) );
  AND2X1 U9414 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[29]), .B(n9038), 
        .Y(n1275) );
  INVX1 U9415 ( .A(n1275), .Y(n7477) );
  AND2X1 U9416 ( .A(recentABools_head_i[3]), .B(ap_CS_fsm[7]), .Y(n1221) );
  INVX1 U9417 ( .A(n1221), .Y(n7478) );
  AND2X1 U9418 ( .A(VbeatFallDelay_new_1_reg_342[10]), .B(n9013), .Y(n2167) );
  INVX1 U9419 ( .A(n2167), .Y(n7479) );
  AND2X1 U9420 ( .A(VbeatFallDelay[12]), .B(n9036), .Y(n1158) );
  INVX1 U9421 ( .A(n1158), .Y(n7480) );
  AND2X1 U9422 ( .A(tmp_5_fu_726_p2[15]), .B(n8993), .Y(n1148) );
  INVX1 U9423 ( .A(n1148), .Y(n7481) );
  AND2X1 U9424 ( .A(VbeatFallDelay_new_1_reg_342[21]), .B(n9013), .Y(n2178) );
  INVX1 U9425 ( .A(n2178), .Y(n7482) );
  AND2X1 U9426 ( .A(VbeatFallDelay[22]), .B(n9035), .Y(n1118) );
  INVX1 U9427 ( .A(n1118), .Y(n7483) );
  AND2X1 U9428 ( .A(VbeatFallDelay_new_1_reg_342[29]), .B(n9013), .Y(n2186) );
  INVX1 U9429 ( .A(n2186), .Y(n7484) );
  AND2X1 U9430 ( .A(tmp_4_fu_716_p2[1]), .B(n8994), .Y(n1075) );
  INVX1 U9431 ( .A(n1075), .Y(n7485) );
  AND2X1 U9432 ( .A(VbeatDelay[4]), .B(n9033), .Y(n1064) );
  INVX1 U9433 ( .A(n1064), .Y(n7486) );
  AND2X1 U9434 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[5]), .Y(n2561) );
  INVX1 U9435 ( .A(n2561), .Y(n7487) );
  AND2X1 U9436 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[14]), .Y(n2552) );
  INVX1 U9437 ( .A(n2552), .Y(n7488) );
  AND2X1 U9438 ( .A(tmp_4_fu_716_p2[20]), .B(n8995), .Y(n1013) );
  INVX1 U9439 ( .A(n1013), .Y(n7489) );
  AND2X1 U9440 ( .A(VbeatDelay[22]), .B(n9032), .Y(n1004) );
  INVX1 U9441 ( .A(n1004), .Y(n7490) );
  AND2X1 U9442 ( .A(VbeatDelay[27]), .B(n9034), .Y(n987) );
  INVX1 U9443 ( .A(n987), .Y(n7491) );
  AND2X1 U9444 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[29]), .Y(n2537) );
  INVX1 U9445 ( .A(n2537), .Y(n7492) );
  BUFX2 U9446 ( .A(n2327), .Y(n7493) );
  AND2X1 U9447 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[18]), .Y(n2478) );
  INVX1 U9448 ( .A(n2478), .Y(n7494) );
  BUFX2 U9449 ( .A(n2314), .Y(n7495) );
  AND2X1 U9450 ( .A(n2273), .B(n9019), .Y(n951) );
  INVX1 U9451 ( .A(n951), .Y(n7496) );
  BUFX2 U9452 ( .A(n2300), .Y(n7497) );
  BUFX2 U9453 ( .A(n2282), .Y(n7498) );
  BUFX2 U9454 ( .A(n2378), .Y(n7499) );
  BUFX2 U9455 ( .A(n2264), .Y(n7500) );
  BUFX2 U9456 ( .A(n2350), .Y(n7501) );
  BUFX2 U9457 ( .A(n2342), .Y(n7502) );
  AND2X1 U9458 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[23]), .B(n970), 
        .Y(n892) );
  INVX1 U9459 ( .A(n892), .Y(n7503) );
  AND2X1 U9460 ( .A(AbeatDelay[3]), .B(n8896), .Y(n781) );
  INVX1 U9461 ( .A(n781), .Y(n7504) );
  AND2X1 U9462 ( .A(AbeatDelay_new_reg_394[5]), .B(n9041), .Y(n2229) );
  INVX1 U9463 ( .A(n2229), .Y(n7505) );
  AND2X1 U9464 ( .A(tmp_3_fu_706_p2[9]), .B(n8996), .Y(n763) );
  INVX1 U9465 ( .A(n763), .Y(n7506) );
  AND2X1 U9466 ( .A(AbeatDelay_new_reg_394[16]), .B(n9041), .Y(n2218) );
  INVX1 U9467 ( .A(n2218), .Y(n7507) );
  AND2X1 U9468 ( .A(AbeatDelay[23]), .B(n10670), .Y(n714) );
  INVX1 U9469 ( .A(n714), .Y(n7508) );
  AND2X1 U9470 ( .A(tmp_3_fu_706_p2[26]), .B(n8997), .Y(n705) );
  INVX1 U9471 ( .A(n705), .Y(n7509) );
  AND2X1 U9472 ( .A(AbeatDelay_new_reg_394[27]), .B(n9041), .Y(n2207) );
  INVX1 U9473 ( .A(n2207), .Y(n7510) );
  AND2X1 U9474 ( .A(AstimDelay[2]), .B(n8896), .Y(n677) );
  INVX1 U9475 ( .A(n677), .Y(n7511) );
  AND2X1 U9476 ( .A(AstimDelay[19]), .B(n8896), .Y(n626) );
  INVX1 U9477 ( .A(n626), .Y(n7512) );
  AND2X1 U9478 ( .A(tmp_6_fu_497_p3[23]), .B(n8966), .Y(n615) );
  INVX1 U9479 ( .A(n615), .Y(n7513) );
  AND2X1 U9480 ( .A(VstimDelay[5]), .B(n10670), .Y(n568) );
  INVX1 U9481 ( .A(n568), .Y(n7514) );
  AND2X1 U9482 ( .A(tmp_7_fu_511_p3[8]), .B(n8965), .Y(n560) );
  INVX1 U9483 ( .A(n560), .Y(n7515) );
  AND2X1 U9484 ( .A(VstimDelay[20]), .B(n8896), .Y(n523) );
  INVX1 U9485 ( .A(n523), .Y(n7516) );
  AND2X1 U9486 ( .A(tmp_7_fu_511_p3[24]), .B(n8963), .Y(n512) );
  INVX1 U9487 ( .A(n512), .Y(n7517) );
  AND2X1 U9488 ( .A(tmp_7_fu_511_p3[27]), .B(n8964), .Y(n503) );
  INVX1 U9489 ( .A(n503), .Y(n7518) );
  AND2X1 U9490 ( .A(VstimDelay[28]), .B(n10670), .Y(n499) );
  INVX1 U9491 ( .A(n499), .Y(n7519) );
  AND2X1 U9492 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[30]), .Y(n2526) );
  INVX1 U9493 ( .A(n2526), .Y(n7520) );
  AND2X1 U9494 ( .A(\Decision_AXILiteS_s_axi_U/n362 ), .B(
        \Decision_AXILiteS_s_axi_U/n351 ), .Y(\Decision_AXILiteS_s_axi_U/n361 ) );
  INVX1 U9495 ( .A(\Decision_AXILiteS_s_axi_U/n361 ), .Y(n7521) );
  AND2X1 U9496 ( .A(a_length[30]), .B(n8116), .Y(
        \Decision_AXILiteS_s_axi_U/n422 ) );
  INVX1 U9497 ( .A(\Decision_AXILiteS_s_axi_U/n422 ), .Y(n7522) );
  AND2X1 U9498 ( .A(\Decision_AXILiteS_s_axi_U/n360 ), .B(n8411), .Y(
        \Decision_AXILiteS_s_axi_U/n464 ) );
  INVX1 U9499 ( .A(\Decision_AXILiteS_s_axi_U/n464 ), .Y(n7523) );
  AND2X1 U9500 ( .A(vthresh[31]), .B(n7865), .Y(
        \Decision_AXILiteS_s_axi_U/n483 ) );
  INVX1 U9501 ( .A(\Decision_AXILiteS_s_axi_U/n483 ), .Y(n7524) );
  AND2X1 U9502 ( .A(s_axi_AXILiteS_AWADDR[3]), .B(n8652), .Y(
        \Decision_AXILiteS_s_axi_U/n638 ) );
  INVX1 U9503 ( .A(\Decision_AXILiteS_s_axi_U/n638 ), .Y(n7525) );
  AND2X1 U9504 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[0]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n379 )
         );
  INVX1 U9505 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n379 ), 
        .Y(n7526) );
  AND2X1 U9506 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[5]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n424 )
         );
  INVX1 U9507 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n424 ), 
        .Y(n7527) );
  AND2X1 U9508 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[11]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n436 )
         );
  INVX1 U9509 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n436 ), 
        .Y(n7528) );
  AND2X1 U9510 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[4]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n456 )
         );
  INVX1 U9511 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n456 ), 
        .Y(n7529) );
  AND2X1 U9512 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[10]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n468 )
         );
  INVX1 U9513 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n468 ), 
        .Y(n7530) );
  AND2X1 U9514 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[3]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n488 )
         );
  INVX1 U9515 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n488 ), 
        .Y(n7531) );
  AND2X1 U9516 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[9]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n500 )
         );
  INVX1 U9517 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n500 ), 
        .Y(n7532) );
  AND2X1 U9518 ( .A(n9467), .B(data_read_reg_1495[2]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n520 )
         );
  INVX1 U9519 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n520 ), 
        .Y(n7533) );
  AND2X1 U9520 ( .A(n9467), .B(data_read_reg_1495[8]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n532 )
         );
  INVX1 U9521 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n532 ), 
        .Y(n7534) );
  AND2X1 U9522 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][6] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n563 )
         );
  INVX1 U9523 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n563 ), 
        .Y(n7535) );
  AND2X1 U9524 ( .A(n9468), .B(data_read_reg_1495[15]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n614 )
         );
  INVX1 U9525 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n614 ), 
        .Y(n7536) );
  AND2X1 U9526 ( .A(n9469), .B(data_read_reg_1495[14]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n646 )
         );
  INVX1 U9527 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n646 ), 
        .Y(n7537) );
  AND2X1 U9528 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][5] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n658 )
         );
  INVX1 U9529 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n658 ), 
        .Y(n7538) );
  AND2X1 U9530 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][4] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n676 )
         );
  INVX1 U9531 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n676 ), 
        .Y(n7539) );
  AND2X1 U9532 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][11] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n701 )
         );
  INVX1 U9533 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n701 ), 
        .Y(n7540) );
  AND2X1 U9534 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][10] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n717 )
         );
  INVX1 U9535 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n717 ), 
        .Y(n7541) );
  AND2X1 U9536 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][9] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n733 )
         );
  INVX1 U9537 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n733 ), 
        .Y(n7542) );
  AND2X1 U9538 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][8] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n749 )
         );
  INVX1 U9539 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n749 ), 
        .Y(n7543) );
  AND2X1 U9540 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][15] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n773 )
         );
  INVX1 U9541 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n773 ), 
        .Y(n7544) );
  AND2X1 U9542 ( .A(n9466), .B(data_read_reg_1495[13]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n802 )
         );
  INVX1 U9543 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n802 ), 
        .Y(n7545) );
  AND2X1 U9544 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][14] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n823 )
         );
  INVX1 U9545 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n823 ), 
        .Y(n7546) );
  AND2X1 U9546 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][1] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n828 )
         );
  INVX1 U9547 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n828 ), 
        .Y(n7547) );
  AND2X1 U9548 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][13] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n840 )
         );
  INVX1 U9549 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n840 ), 
        .Y(n7548) );
  AND2X1 U9550 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][0] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n844 )
         );
  INVX1 U9551 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n844 ), 
        .Y(n7549) );
  AND2X1 U9552 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][12] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n856 )
         );
  INVX1 U9553 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n856 ), 
        .Y(n7550) );
  AND2X1 U9554 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[12]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n886 )
         );
  INVX1 U9555 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n886 ), 
        .Y(n7551) );
  BUFX2 U9556 ( .A(n11814), .Y(n7552) );
  AND2X1 U9557 ( .A(sum_reg_308[30]), .B(n8929), .Y(n2578) );
  INVX1 U9558 ( .A(n2578), .Y(n7553) );
  AND2X1 U9559 ( .A(tmp_29_i_fu_752_p2[14]), .B(n8920), .Y(n3179) );
  INVX1 U9560 ( .A(n3179), .Y(n7554) );
  AND2X1 U9561 ( .A(tmp_29_i1_fu_1065_p2[14]), .B(n8922), .Y(n3231) );
  INVX1 U9562 ( .A(n3231), .Y(n7555) );
  AND2X1 U9563 ( .A(tmp_29_i_fu_752_p2[4]), .B(n8920), .Y(n3158) );
  INVX1 U9564 ( .A(n3158), .Y(n7556) );
  AND2X1 U9565 ( .A(tmp_29_i1_fu_1065_p2[4]), .B(n8922), .Y(n3210) );
  INVX1 U9566 ( .A(n3210), .Y(n7557) );
  AND2X1 U9567 ( .A(CircularBuffer_len_write_assig_fu_817_p2[11]), .B(n8894), 
        .Y(n1587) );
  INVX1 U9568 ( .A(n1587), .Y(n7558) );
  AND2X1 U9569 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[11]), .B(n8891), .Y(n911) );
  INVX1 U9570 ( .A(n911), .Y(n7559) );
  AND2X1 U9571 ( .A(sum_1_reg_376[6]), .B(n8930), .Y(n2432) );
  INVX1 U9572 ( .A(n2432), .Y(n7560) );
  AND2X1 U9573 ( .A(sum_reg_308[9]), .B(n8929), .Y(n2662) );
  INVX1 U9574 ( .A(n2662), .Y(n7561) );
  AND2X1 U9575 ( .A(sum_1_reg_376[21]), .B(n8930), .Y(n2492) );
  INVX1 U9576 ( .A(n2492), .Y(n7562) );
  INVX1 U9577 ( .A(n3861), .Y(n7563) );
  AND2X1 U9578 ( .A(CircularBuffer_head_i_read_ass_reg_1624[4]), .B(n9008), 
        .Y(n1709) );
  INVX1 U9579 ( .A(n1709), .Y(n7564) );
  INVX1 U9580 ( .A(n3656), .Y(n7565) );
  AND2X1 U9581 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[3]), .B(n9037), 
        .Y(n1224) );
  INVX1 U9582 ( .A(n1224), .Y(n7566) );
  BUFX2 U9583 ( .A(n12189), .Y(n7567) );
  AND2X1 U9584 ( .A(v_thresh[18]), .B(n9540), .Y(n12187) );
  INVX1 U9585 ( .A(n12187), .Y(n7568) );
  BUFX2 U9586 ( .A(n11556), .Y(n7569) );
  AND2X1 U9587 ( .A(a_thresh[18]), .B(n9490), .Y(n11554) );
  INVX1 U9588 ( .A(n11554), .Y(n7570) );
  INVX1 U9589 ( .A(n4618), .Y(n7571) );
  AND2X1 U9590 ( .A(ACaptureThresh_loc_reg_288[16]), .B(n8968), .Y(n3030) );
  INVX1 U9591 ( .A(n3030), .Y(n7572) );
  BUFX2 U9592 ( .A(n3029), .Y(n7573) );
  INVX1 U9593 ( .A(n4603), .Y(n7574) );
  AND2X1 U9594 ( .A(ACaptureThresh_loc_reg_288[31]), .B(n8971), .Y(n3000) );
  INVX1 U9595 ( .A(n3000), .Y(n7575) );
  BUFX2 U9596 ( .A(n2999), .Y(n7576) );
  INVX1 U9597 ( .A(n4555), .Y(n7577) );
  AND2X1 U9598 ( .A(VCaptureThresh_loc_reg_298[15]), .B(n8970), .Y(n2904) );
  INVX1 U9599 ( .A(n2904), .Y(n7578) );
  BUFX2 U9600 ( .A(n2903), .Y(n7579) );
  INVX1 U9601 ( .A(n4542), .Y(n7580) );
  AND2X1 U9602 ( .A(VCaptureThresh_loc_reg_298[28]), .B(n8969), .Y(n2878) );
  INVX1 U9603 ( .A(n2878), .Y(n7581) );
  BUFX2 U9604 ( .A(n2877), .Y(n7582) );
  INVX1 U9605 ( .A(n12252), .Y(n7583) );
  BUFX2 U9606 ( .A(n12251), .Y(n7584) );
  INVX1 U9607 ( .A(n11619), .Y(n7585) );
  BUFX2 U9608 ( .A(n11618), .Y(n7586) );
  INVX1 U9609 ( .A(n11916), .Y(n7587) );
  BUFX2 U9610 ( .A(n11915), .Y(n7588) );
  OR2X1 U9611 ( .A(VbeatFallDelay_new_1_reg_342[14]), .B(
        VbeatFallDelay_new_1_reg_342[13]), .Y(n11914) );
  INVX1 U9612 ( .A(n11914), .Y(n7589) );
  OR2X1 U9613 ( .A(p_tmp_i_reg_1556[20]), .B(p_tmp_i_reg_1556[19]), .Y(n11245)
         );
  INVX1 U9614 ( .A(n11245), .Y(n7590) );
  BUFX2 U9615 ( .A(n11093), .Y(n7591) );
  AND2X1 U9616 ( .A(VbeatDelay_new_1_reg_326[9]), .B(n10697), .Y(n11092) );
  INVX1 U9617 ( .A(n11092), .Y(n7592) );
  AND2X1 U9618 ( .A(n10274), .B(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n9 ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n8 ) );
  INVX1 U9619 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n8 ), 
        .Y(n7593) );
  BUFX2 U9620 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n7 ), 
        .Y(n7594) );
  BUFX2 U9621 ( .A(n11167), .Y(n7595) );
  BUFX2 U9622 ( .A(n11157), .Y(n7596) );
  BUFX2 U9623 ( .A(n11890), .Y(n7597) );
  BUFX2 U9624 ( .A(n11888), .Y(n7598) );
  AND2X1 U9625 ( .A(n9909), .B(n9908), .Y(n1689) );
  INVX1 U9626 ( .A(n1689), .Y(n7599) );
  AND2X1 U9627 ( .A(n10093), .B(n10094), .Y(n1486) );
  INVX1 U9628 ( .A(n1486), .Y(n7600) );
  AND2X1 U9629 ( .A(n10588), .B(n10589), .Y(n851) );
  INVX1 U9630 ( .A(n851), .Y(n7601) );
  AND2X1 U9631 ( .A(n10705), .B(n10707), .Y(n269) );
  INVX1 U9632 ( .A(n269), .Y(n7602) );
  AND2X1 U9633 ( .A(n10132), .B(n10133), .Y(n3204) );
  INVX1 U9634 ( .A(n3204), .Y(n7603) );
  AND2X1 U9635 ( .A(n10627), .B(n10628), .Y(n3256) );
  INVX1 U9636 ( .A(n3256), .Y(n7604) );
  AND2X1 U9637 ( .A(n9906), .B(n9905), .Y(n2070) );
  INVX1 U9638 ( .A(n2070), .Y(n7605) );
  BUFX2 U9639 ( .A(n1521), .Y(n7606) );
  OR2X1 U9640 ( .A(CircularBuffer_len_write_assig_reg_1634[2]), .B(
        CircularBuffer_len_write_assig_reg_1634[29]), .Y(n1528) );
  INVX1 U9641 ( .A(n1528), .Y(n7607) );
  BUFX2 U9642 ( .A(n799), .Y(n7608) );
  OR2X1 U9643 ( .A(CircularBuffer_len_write_assig_2_reg_1729[2]), .B(
        CircularBuffer_len_write_assig_2_reg_1729[29]), .Y(n806) );
  INVX1 U9644 ( .A(n806), .Y(n7609) );
  AND2X1 U9645 ( .A(n10463), .B(n10466), .Y(n330) );
  INVX1 U9646 ( .A(n330), .Y(n7610) );
  BUFX2 U9647 ( .A(n328), .Y(n7611) );
  BUFX2 U9648 ( .A(n329), .Y(n7612) );
  AND2X1 U9649 ( .A(n9840), .B(n9841), .Y(n2034) );
  INVX1 U9650 ( .A(n2034), .Y(n7613) );
  AND2X1 U9651 ( .A(n9838), .B(n9839), .Y(n2035) );
  INVX1 U9652 ( .A(n2035), .Y(n7614) );
  BUFX2 U9653 ( .A(n2033), .Y(n7615) );
  AND2X1 U9654 ( .A(n11233), .B(n7861), .Y(n11234) );
  INVX1 U9655 ( .A(n11234), .Y(n7616) );
  AND2X1 U9656 ( .A(n11203), .B(n7862), .Y(n11204) );
  INVX1 U9657 ( .A(n11204), .Y(n7617) );
  AND2X1 U9658 ( .A(n11231), .B(n8111), .Y(n11232) );
  INVX1 U9659 ( .A(n11232), .Y(n7618) );
  AND2X1 U9660 ( .A(n11201), .B(n8112), .Y(n11202) );
  INVX1 U9661 ( .A(n11202), .Y(n7619) );
  AND2X1 U9662 ( .A(n11209), .B(n8113), .Y(n11210) );
  INVX1 U9663 ( .A(n11210), .Y(n7620) );
  AND2X1 U9664 ( .A(n11179), .B(n8114), .Y(n11180) );
  INVX1 U9665 ( .A(n11180), .Y(n7621) );
  AND2X1 U9666 ( .A(recentdatapoints_len_load_op_fu_556_p2[11]), .B(n8972), 
        .Y(n1833) );
  INVX1 U9667 ( .A(n1833), .Y(n7622) );
  AND2X1 U9668 ( .A(recentdatapoints_len_load_op_fu_556_p2[24]), .B(n8972), 
        .Y(n1849) );
  INVX1 U9669 ( .A(n1849), .Y(n7623) );
  AND2X1 U9670 ( .A(recentdatapoints_len_load_op_fu_556_p2[28]), .B(n8972), 
        .Y(n1855) );
  INVX1 U9671 ( .A(n1855), .Y(n7624) );
  AND2X1 U9672 ( .A(ap_rst_n), .B(n8388), .Y(\Decision_AXILiteS_s_axi_U/n600 )
         );
  INVX1 U9673 ( .A(\Decision_AXILiteS_s_axi_U/n600 ), .Y(n7625) );
  BUFX2 U9674 ( .A(n1865), .Y(n7626) );
  AND2X1 U9675 ( .A(n9935), .B(tmp_33_i_fu_786_p2[3]), .Y(n1703) );
  INVX1 U9676 ( .A(n1703), .Y(n7627) );
  AND2X1 U9677 ( .A(n10243), .B(tmp_33_i1_fu_1099_p2[4]), .Y(n1228) );
  INVX1 U9678 ( .A(n1228), .Y(n7628) );
  BUFX2 U9679 ( .A(n11602), .Y(n7629) );
  BUFX2 U9680 ( .A(n2196), .Y(n7630) );
  OR2X1 U9681 ( .A(i_5_fu_854_p2[3]), .B(n8641), .Y(n8848) );
  BUFX2 U9682 ( .A(\Decision_AXILiteS_s_axi_U/n615 ), .Y(n7631) );
  OR2X1 U9683 ( .A(n9677), .B(n2776), .Y(n12116) );
  INVX1 U9684 ( .A(n12116), .Y(n7632) );
  OR2X1 U9685 ( .A(n9573), .B(n2283), .Y(n11652) );
  INVX1 U9686 ( .A(n11652), .Y(n7633) );
  BUFX2 U9687 ( .A(n11367), .Y(n7634) );
  BUFX2 U9688 ( .A(n11368), .Y(n7635) );
  BUFX2 U9689 ( .A(n11419), .Y(n7636) );
  BUFX2 U9690 ( .A(n11420), .Y(n7637) );
  AND2X1 U9691 ( .A(recentdatapoints_data_q0[3]), .B(n8869), .Y(n412) );
  INVX1 U9692 ( .A(n412), .Y(n7638) );
  AND2X1 U9693 ( .A(recentdatapoints_data_q0[13]), .B(n8868), .Y(n421) );
  INVX1 U9694 ( .A(n421), .Y(n7639) );
  AND2X1 U9695 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[4]), 
        .Y(n452) );
  INVX1 U9696 ( .A(n452), .Y(n7640) );
  AND2X1 U9697 ( .A(CircularBuffer_len_read_assign_fu_772_p2[13]), .B(n3151), 
        .Y(n2768) );
  INVX1 U9698 ( .A(n2768), .Y(n7641) );
  AND2X1 U9699 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[13]), .B(n3149), .Y(n2275) );
  INVX1 U9700 ( .A(n2275), .Y(n7642) );
  AND2X1 U9701 ( .A(CircularBuffer_len_read_assign_fu_772_p2[6]), .B(n3151), 
        .Y(n2782) );
  INVX1 U9702 ( .A(n2782), .Y(n7643) );
  AND2X1 U9703 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[6]), .B(n3149), 
        .Y(n2289) );
  INVX1 U9704 ( .A(n2289), .Y(n7644) );
  AND2X1 U9705 ( .A(CircularBuffer_len_read_assign_fu_772_p2[27]), .B(n8919), 
        .Y(n2740) );
  INVX1 U9706 ( .A(n2740), .Y(n7645) );
  AND2X1 U9707 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[27]), .B(n8921), .Y(n2247) );
  INVX1 U9708 ( .A(n2247), .Y(n7646) );
  AND2X1 U9709 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n71 ), .B(recentVBools_data_address0[0]), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n46 ) );
  INVX1 U9710 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n46 ), 
        .Y(n7647) );
  AND2X1 U9711 ( .A(recentVBools_data_address0[1]), .B(n8413), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n71 ) );
  INVX1 U9712 ( .A(recentABools_data_address0[2]), .Y(n7648) );
  BUFX2 U9713 ( .A(n390), .Y(n7649) );
  BUFX2 U9714 ( .A(n391), .Y(n7650) );
  AND2X1 U9715 ( .A(\Decision_AXILiteS_s_axi_U/n533 ), .B(
        \Decision_AXILiteS_s_axi_U/n384 ), .Y(\Decision_AXILiteS_s_axi_U/n525 ) );
  INVX1 U9716 ( .A(\Decision_AXILiteS_s_axi_U/n525 ), .Y(n7651) );
  AND2X1 U9717 ( .A(\Decision_AXILiteS_s_axi_U/n385 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n373 ) );
  INVX1 U9718 ( .A(\Decision_AXILiteS_s_axi_U/n373 ), .Y(n7652) );
  AND2X1 U9719 ( .A(n10060), .B(\tmp_12_reg_1694[0] ), .Y(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n35 ) );
  INVX1 U9720 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n35 ), 
        .Y(n7653) );
  BUFX2 U9721 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n36 ), 
        .Y(n7654) );
  AND2X1 U9722 ( .A(\Decision_AXILiteS_s_axi_U/n397 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n430 ) );
  INVX1 U9723 ( .A(\Decision_AXILiteS_s_axi_U/n430 ), .Y(n7655) );
  AND2X1 U9724 ( .A(\Decision_AXILiteS_s_axi_U/n353 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n503 ) );
  INVX1 U9725 ( .A(\Decision_AXILiteS_s_axi_U/n503 ), .Y(n7656) );
  AND2X1 U9726 ( .A(a_length[0]), .B(n8951), .Y(n3126) );
  INVX1 U9727 ( .A(n3126), .Y(n7657) );
  AND2X1 U9728 ( .A(a_length[12]), .B(n8952), .Y(n3102) );
  INVX1 U9729 ( .A(n3102), .Y(n7658) );
  AND2X1 U9730 ( .A(v_length[6]), .B(n8954), .Y(n2986) );
  INVX1 U9731 ( .A(n2986), .Y(n7659) );
  AND2X1 U9732 ( .A(v_length[22]), .B(n8955), .Y(n2954) );
  INVX1 U9733 ( .A(n2954), .Y(n7660) );
  AND2X1 U9734 ( .A(a_flip[0]), .B(n8953), .Y(n2869) );
  INVX1 U9735 ( .A(n2869), .Y(n7661) );
  AND2X1 U9736 ( .A(recentdatapoints_head_i[31]), .B(n8979), .Y(n1952) );
  INVX1 U9737 ( .A(n1952), .Y(n7662) );
  AND2X1 U9738 ( .A(p_tmp_i_reg_1556[19]), .B(n8980), .Y(n1900) );
  INVX1 U9739 ( .A(n1900), .Y(n7663) );
  AND2X1 U9740 ( .A(p_tmp_i_reg_1556[7]), .B(n8980), .Y(n1876) );
  INVX1 U9741 ( .A(n1876), .Y(n7664) );
  AND2X1 U9742 ( .A(CircularBuffer_head_i_read_ass_reg_1624[18]), .B(n9010), 
        .Y(n1751) );
  INVX1 U9743 ( .A(n1751), .Y(n7665) );
  AND2X1 U9744 ( .A(CircularBuffer_head_i_read_ass_reg_1624[26]), .B(n9009), 
        .Y(n1727) );
  INVX1 U9745 ( .A(n1727), .Y(n7666) );
  AND2X1 U9746 ( .A(ap_CS_fsm[2]), .B(recentVBools_head_i[4]), .Y(n1706) );
  INVX1 U9747 ( .A(n1706), .Y(n7667) );
  BUFX2 U9748 ( .A(n2815), .Y(n7668) );
  AND2X1 U9749 ( .A(CircularBuffer_len_write_assig_fu_817_p2[8]), .B(n8894), 
        .Y(n1591) );
  INVX1 U9750 ( .A(n1591), .Y(n7669) );
  BUFX2 U9751 ( .A(n2797), .Y(n7670) );
  BUFX2 U9752 ( .A(n2795), .Y(n7671) );
  AND2X1 U9753 ( .A(CircularBuffer_sum_read_assign_reg_1610[28]), .B(n9006), 
        .Y(n1410) );
  INVX1 U9754 ( .A(n1410), .Y(n7672) );
  AND2X1 U9755 ( .A(CircularBuffer_sum_read_assign_reg_1610[31]), .B(n9007), 
        .Y(n1404) );
  INVX1 U9756 ( .A(n1404), .Y(n7673) );
  BUFX2 U9757 ( .A(n2729), .Y(n7674) );
  AND2X1 U9758 ( .A(n9012), .B(sum_phi_fu_311_p4[15]), .Y(n2636) );
  INVX1 U9759 ( .A(n2636), .Y(n7675) );
  BUFX2 U9760 ( .A(n2716), .Y(n7676) );
  BUFX2 U9761 ( .A(n2703), .Y(n7677) );
  AND2X1 U9762 ( .A(recentABools_head_i[12]), .B(n9040), .Y(n1314) );
  INVX1 U9763 ( .A(n1314), .Y(n7678) );
  AND2X1 U9764 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[19]), .B(n9039), 
        .Y(n1301) );
  INVX1 U9765 ( .A(n1301), .Y(n7679) );
  AND2X1 U9766 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[25]), .B(n9038), 
        .Y(n1285) );
  INVX1 U9767 ( .A(n1285), .Y(n7680) );
  AND2X1 U9768 ( .A(recentABools_head_i[2]), .B(ap_CS_fsm[7]), .Y(n1216) );
  INVX1 U9769 ( .A(n1216), .Y(n7681) );
  AND2X1 U9770 ( .A(n10365), .B(n8992), .Y(n1206) );
  INVX1 U9771 ( .A(n1206), .Y(n7682) );
  AND2X1 U9772 ( .A(VbeatFallDelay_new_1_reg_342[11]), .B(n9013), .Y(n2168) );
  INVX1 U9773 ( .A(n2168), .Y(n7683) );
  AND2X1 U9774 ( .A(VbeatFallDelay[13]), .B(n9036), .Y(n1154) );
  INVX1 U9775 ( .A(n1154), .Y(n7684) );
  AND2X1 U9776 ( .A(tmp_5_fu_726_p2[16]), .B(n8993), .Y(n1144) );
  INVX1 U9777 ( .A(n1144), .Y(n7685) );
  AND2X1 U9778 ( .A(VbeatFallDelay_new_1_reg_342[22]), .B(n9013), .Y(n2179) );
  INVX1 U9779 ( .A(n2179), .Y(n7686) );
  AND2X1 U9780 ( .A(VbeatFallDelay_new_1_reg_342[30]), .B(n9013), .Y(n2187) );
  INVX1 U9781 ( .A(n2187), .Y(n7687) );
  AND2X1 U9782 ( .A(tmp_4_fu_716_p2[2]), .B(n8994), .Y(n1071) );
  INVX1 U9783 ( .A(n1071), .Y(n7688) );
  AND2X1 U9784 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[3]), .Y(n2563) );
  INVX1 U9785 ( .A(n2563), .Y(n7689) );
  AND2X1 U9786 ( .A(VbeatDelay[7]), .B(n9033), .Y(n1054) );
  INVX1 U9787 ( .A(n1054), .Y(n7690) );
  AND2X1 U9788 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[15]), .Y(n2551) );
  INVX1 U9789 ( .A(n2551), .Y(n7691) );
  AND2X1 U9790 ( .A(tmp_4_fu_716_p2[21]), .B(n8995), .Y(n1009) );
  INVX1 U9791 ( .A(n1009), .Y(n7692) );
  AND2X1 U9792 ( .A(VbeatDelay[23]), .B(n9032), .Y(n1001) );
  INVX1 U9793 ( .A(n1001), .Y(n7693) );
  AND2X1 U9794 ( .A(VbeatDelay[28]), .B(n9034), .Y(n983) );
  INVX1 U9795 ( .A(n983), .Y(n7694) );
  AND2X1 U9796 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[31]), .Y(n2534) );
  INVX1 U9797 ( .A(n2534), .Y(n7695) );
  BUFX2 U9798 ( .A(n2326), .Y(n7696) );
  AND2X1 U9799 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[19]), .Y(n2482) );
  INVX1 U9800 ( .A(n2482), .Y(n7697) );
  BUFX2 U9801 ( .A(n2312), .Y(n7698) );
  AND2X1 U9802 ( .A(n9017), .B(CircularBuffer_len_read_assign_3_fu_1091_p3[2]), 
        .Y(n967) );
  INVX1 U9803 ( .A(n967), .Y(n7699) );
  AND2X1 U9804 ( .A(n2238), .B(n9019), .Y(n928) );
  INVX1 U9805 ( .A(n928), .Y(n7700) );
  BUFX2 U9806 ( .A(n2376), .Y(n7701) );
  BUFX2 U9807 ( .A(n2348), .Y(n7702) );
  AND2X1 U9808 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[8]), .B(n8891), 
        .Y(n915) );
  INVX1 U9809 ( .A(n915), .Y(n7703) );
  BUFX2 U9810 ( .A(n2302), .Y(n7704) );
  AND2X1 U9811 ( .A(AbeatDelay_new_reg_394[4]), .B(n9041), .Y(n2230) );
  INVX1 U9812 ( .A(n2230), .Y(n7705) );
  AND2X1 U9813 ( .A(tmp_3_fu_706_p2[10]), .B(n8996), .Y(n760) );
  INVX1 U9814 ( .A(n760), .Y(n7706) );
  AND2X1 U9815 ( .A(AbeatDelay_new_reg_394[17]), .B(n9041), .Y(n2217) );
  INVX1 U9816 ( .A(n2217), .Y(n7707) );
  AND2X1 U9817 ( .A(AbeatDelay[22]), .B(n10670), .Y(n717) );
  INVX1 U9818 ( .A(n717), .Y(n7708) );
  AND2X1 U9819 ( .A(tmp_3_fu_706_p2[23]), .B(n8997), .Y(n716) );
  INVX1 U9820 ( .A(n716), .Y(n7709) );
  AND2X1 U9821 ( .A(AbeatDelay_new_reg_394[28]), .B(n9041), .Y(n2206) );
  INVX1 U9822 ( .A(n2206), .Y(n7710) );
  AND2X1 U9823 ( .A(tmp_3_fu_706_p2[30]), .B(ap_CS_fsm[4]), .Y(n691) );
  INVX1 U9824 ( .A(n691), .Y(n7711) );
  AND2X1 U9825 ( .A(AstimDelay[3]), .B(n10670), .Y(n674) );
  INVX1 U9826 ( .A(n674), .Y(n7712) );
  AND2X1 U9827 ( .A(tmp_6_fu_497_p3[6]), .B(n8967), .Y(n666) );
  INVX1 U9828 ( .A(n666), .Y(n7713) );
  AND2X1 U9829 ( .A(AstimDelay[20]), .B(n8896), .Y(n623) );
  INVX1 U9830 ( .A(n623), .Y(n7714) );
  AND2X1 U9831 ( .A(tmp_6_fu_497_p3[24]), .B(n8966), .Y(n612) );
  INVX1 U9832 ( .A(n612), .Y(n7715) );
  AND2X1 U9833 ( .A(VstimDelay[6]), .B(n8896), .Y(n565) );
  INVX1 U9834 ( .A(n565), .Y(n7716) );
  AND2X1 U9835 ( .A(VstimDelay[21]), .B(n8896), .Y(n520) );
  INVX1 U9836 ( .A(n520), .Y(n7717) );
  AND2X1 U9837 ( .A(tmp_7_fu_511_p3[28]), .B(n8964), .Y(n500) );
  INVX1 U9838 ( .A(n500), .Y(n7718) );
  AND2X1 U9839 ( .A(VstimDelay[29]), .B(n10670), .Y(n496) );
  INVX1 U9840 ( .A(n496), .Y(n7719) );
  AND2X1 U9841 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[31]), .B(n9035), 
        .Y(n483) );
  INVX1 U9842 ( .A(n483), .Y(n7720) );
  AND2X1 U9843 ( .A(\Decision_AXILiteS_s_axi_U/n356 ), .B(
        \Decision_AXILiteS_s_axi_U/n351 ), .Y(\Decision_AXILiteS_s_axi_U/n355 ) );
  INVX1 U9844 ( .A(\Decision_AXILiteS_s_axi_U/n355 ), .Y(n7721) );
  AND2X1 U9845 ( .A(\Decision_AXILiteS_s_axi_U/n358 ), .B(n8411), .Y(
        \Decision_AXILiteS_s_axi_U/n463 ) );
  INVX1 U9846 ( .A(\Decision_AXILiteS_s_axi_U/n463 ), .Y(n7722) );
  AND2X1 U9847 ( .A(s_axi_AXILiteS_AWADDR[4]), .B(n8652), .Y(
        \Decision_AXILiteS_s_axi_U/n639 ) );
  INVX1 U9848 ( .A(\Decision_AXILiteS_s_axi_U/n639 ), .Y(n7723) );
  AND2X1 U9849 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[1]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n381 )
         );
  INVX1 U9850 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n381 ), 
        .Y(n7724) );
  AND2X1 U9851 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[4]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n422 )
         );
  INVX1 U9852 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n422 ), 
        .Y(n7725) );
  AND2X1 U9853 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[10]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n434 )
         );
  INVX1 U9854 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n434 ), 
        .Y(n7726) );
  AND2X1 U9855 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[5]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n458 )
         );
  INVX1 U9856 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n458 ), 
        .Y(n7727) );
  AND2X1 U9857 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[11]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n470 )
         );
  INVX1 U9858 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n470 ), 
        .Y(n7728) );
  AND2X1 U9859 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[2]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n486 )
         );
  INVX1 U9860 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n486 ), 
        .Y(n7729) );
  AND2X1 U9861 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[8]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n498 )
         );
  INVX1 U9862 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n498 ), 
        .Y(n7730) );
  AND2X1 U9863 ( .A(n9467), .B(data_read_reg_1495[3]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n522 )
         );
  INVX1 U9864 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n522 ), 
        .Y(n7731) );
  AND2X1 U9865 ( .A(n9467), .B(data_read_reg_1495[9]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n534 )
         );
  INVX1 U9866 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n534 ), 
        .Y(n7732) );
  AND2X1 U9867 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][7] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n565 )
         );
  INVX1 U9868 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n565 ), 
        .Y(n7733) );
  AND2X1 U9869 ( .A(n9468), .B(data_read_reg_1495[14]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n612 )
         );
  INVX1 U9870 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n612 ), 
        .Y(n7734) );
  AND2X1 U9871 ( .A(n9469), .B(data_read_reg_1495[15]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n648 )
         );
  INVX1 U9872 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n648 ), 
        .Y(n7735) );
  AND2X1 U9873 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][4] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n657 )
         );
  INVX1 U9874 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n657 ), 
        .Y(n7736) );
  AND2X1 U9875 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][5] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n677 )
         );
  INVX1 U9876 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n677 ), 
        .Y(n7737) );
  AND2X1 U9877 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][10] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n700 )
         );
  INVX1 U9878 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n700 ), 
        .Y(n7738) );
  AND2X1 U9879 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][11] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n718 )
         );
  INVX1 U9880 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n718 ), 
        .Y(n7739) );
  AND2X1 U9881 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][8] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n732 )
         );
  INVX1 U9882 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n732 ), 
        .Y(n7740) );
  AND2X1 U9883 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][9] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n750 )
         );
  INVX1 U9884 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n750 ), 
        .Y(n7741) );
  AND2X1 U9885 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][14] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n772 )
         );
  INVX1 U9886 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n772 ), 
        .Y(n7742) );
  AND2X1 U9887 ( .A(n9466), .B(data_read_reg_1495[12]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n800 )
         );
  INVX1 U9888 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n800 ), 
        .Y(n7743) );
  AND2X1 U9889 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][15] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n824 )
         );
  INVX1 U9890 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n824 ), 
        .Y(n7744) );
  AND2X1 U9891 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][0] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n827 )
         );
  INVX1 U9892 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n827 ), 
        .Y(n7745) );
  AND2X1 U9893 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][12] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n839 )
         );
  INVX1 U9894 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n839 ), 
        .Y(n7746) );
  AND2X1 U9895 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][1] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n845 )
         );
  INVX1 U9896 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n845 ), 
        .Y(n7747) );
  AND2X1 U9897 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][13] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n857 )
         );
  INVX1 U9898 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n857 ), 
        .Y(n7748) );
  AND2X1 U9899 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[13]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n888 )
         );
  INVX1 U9900 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n888 ), 
        .Y(n7749) );
  AND2X1 U9901 ( .A(sum_reg_308[27]), .B(n8929), .Y(n2590) );
  INVX1 U9902 ( .A(n2590), .Y(n7750) );
  AND2X1 U9903 ( .A(tmp_6_fu_497_p3[31]), .B(n8965), .Y(n591) );
  INVX1 U9904 ( .A(n591), .Y(n7751) );
  AND2X1 U9905 ( .A(n471), .B(n439), .Y(n472) );
  INVX1 U9906 ( .A(n472), .Y(n7752) );
  AND2X1 U9907 ( .A(tmp_29_i_fu_752_p2[13]), .B(n8920), .Y(n3180) );
  INVX1 U9908 ( .A(n3180), .Y(n7753) );
  AND2X1 U9909 ( .A(tmp_29_i1_fu_1065_p2[13]), .B(n8922), .Y(n3232) );
  INVX1 U9910 ( .A(n3232), .Y(n7754) );
  AND2X1 U9911 ( .A(tmp_29_i_fu_752_p2[3]), .B(n8920), .Y(n3159) );
  INVX1 U9912 ( .A(n3159), .Y(n7755) );
  AND2X1 U9913 ( .A(tmp_29_i1_fu_1065_p2[3]), .B(n8922), .Y(n3211) );
  INVX1 U9914 ( .A(n3211), .Y(n7756) );
  AND2X1 U9915 ( .A(N502), .B(ap_CS_fsm[12]), .Y(n590) );
  INVX1 U9916 ( .A(n590), .Y(n7757) );
  AND2X1 U9917 ( .A(sum_1_reg_376[5]), .B(n8930), .Y(n2428) );
  INVX1 U9918 ( .A(n2428), .Y(n7758) );
  AND2X1 U9919 ( .A(sum_reg_308[6]), .B(n8929), .Y(n2674) );
  INVX1 U9920 ( .A(n2674), .Y(n7759) );
  AND2X1 U9921 ( .A(sum_1_reg_376[18]), .B(n8930), .Y(n2480) );
  INVX1 U9922 ( .A(n2480), .Y(n7760) );
  INVX1 U9923 ( .A(n3857), .Y(n7761) );
  AND2X1 U9924 ( .A(CircularBuffer_head_i_read_ass_reg_1624[2]), .B(n9008), 
        .Y(n1702) );
  INVX1 U9925 ( .A(n1702), .Y(n7762) );
  INVX1 U9926 ( .A(n3653), .Y(n7763) );
  AND2X1 U9927 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[2]), .B(n9037), 
        .Y(n1219) );
  INVX1 U9928 ( .A(n1219), .Y(n7764) );
  INVX1 U9929 ( .A(n4617), .Y(n7765) );
  AND2X1 U9930 ( .A(ACaptureThresh_loc_reg_288[17]), .B(n8969), .Y(n3028) );
  INVX1 U9931 ( .A(n3028), .Y(n7766) );
  BUFX2 U9932 ( .A(n3027), .Y(n7767) );
  INVX1 U9933 ( .A(n4570), .Y(n7768) );
  AND2X1 U9934 ( .A(VCaptureThresh_loc_reg_298[0]), .B(n8971), .Y(n2934) );
  INVX1 U9935 ( .A(n2934), .Y(n7769) );
  BUFX2 U9936 ( .A(n2933), .Y(n7770) );
  INVX1 U9937 ( .A(n4557), .Y(n7771) );
  AND2X1 U9938 ( .A(VCaptureThresh_loc_reg_298[13]), .B(n8970), .Y(n2908) );
  INVX1 U9939 ( .A(n2908), .Y(n7772) );
  BUFX2 U9940 ( .A(n2907), .Y(n7773) );
  INVX1 U9941 ( .A(n4541), .Y(n7774) );
  AND2X1 U9942 ( .A(VCaptureThresh_loc_reg_298[29]), .B(n8969), .Y(n2876) );
  INVX1 U9943 ( .A(n2876), .Y(n7775) );
  BUFX2 U9944 ( .A(n2875), .Y(n7776) );
  BUFX2 U9945 ( .A(n12190), .Y(n7777) );
  AND2X1 U9946 ( .A(v_thresh[17]), .B(n9540), .Y(n12185) );
  INVX1 U9947 ( .A(n12185), .Y(n7778) );
  BUFX2 U9948 ( .A(n11557), .Y(n7779) );
  AND2X1 U9949 ( .A(a_thresh[17]), .B(n9490), .Y(n11552) );
  INVX1 U9950 ( .A(n11552), .Y(n7780) );
  OR2X1 U9951 ( .A(n8087), .B(v_thresh[30]), .Y(n12249) );
  INVX1 U9952 ( .A(n12249), .Y(n7781) );
  OR2X1 U9953 ( .A(n8088), .B(a_thresh[30]), .Y(n11616) );
  INVX1 U9954 ( .A(n11616), .Y(n7782) );
  BUFX2 U9955 ( .A(n11925), .Y(n7783) );
  AND2X1 U9956 ( .A(tmp_6_reg_1538[9]), .B(n9573), .Y(n11924) );
  INVX1 U9957 ( .A(n11924), .Y(n7784) );
  BUFX2 U9958 ( .A(n12014), .Y(n7785) );
  AND2X1 U9959 ( .A(tmp_7_reg_1544[9]), .B(n9677), .Y(n12013) );
  INVX1 U9960 ( .A(n12013), .Y(n7786) );
  BUFX2 U9961 ( .A(n11817), .Y(n7787) );
  AND2X1 U9962 ( .A(VbeatDelay_new_1_reg_326[9]), .B(n10390), .Y(n11816) );
  INVX1 U9963 ( .A(n11816), .Y(n7788) );
  AND2X1 U9964 ( .A(VbeatDelay_new_1_reg_326[29]), .B(n10737), .Y(n11145) );
  INVX1 U9965 ( .A(n11145), .Y(n7789) );
  AND2X1 U9966 ( .A(n11902), .B(n11901), .Y(n11907) );
  INVX1 U9967 ( .A(n11907), .Y(n7790) );
  BUFX2 U9968 ( .A(n11906), .Y(n7791) );
  BUFX2 U9969 ( .A(n11844), .Y(n7792) );
  BUFX2 U9970 ( .A(n11891), .Y(n7793) );
  BUFX2 U9971 ( .A(n11881), .Y(n7794) );
  OR2X1 U9972 ( .A(n9995), .B(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n140 ), .Y(
        \recentVBools_data_U/Decision_recentVBools_data_ram_U/n144 ) );
  INVX1 U9973 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n144 ), .Y(n7795) );
  BUFX2 U9974 ( .A(n12088), .Y(n7796) );
  BUFX2 U9975 ( .A(n12078), .Y(n7797) );
  AND2X1 U9976 ( .A(n9012), .B(n9859), .Y(n1668) );
  INVX1 U9977 ( .A(n1668), .Y(n7798) );
  AND2X1 U9978 ( .A(n10080), .B(n10108), .Y(n1505) );
  INVX1 U9979 ( .A(n1505), .Y(n7799) );
  AND2X1 U9980 ( .A(n9862), .B(n9861), .Y(n1950) );
  INVX1 U9981 ( .A(n1950), .Y(n7800) );
  AND2X1 U9982 ( .A(n10729), .B(n10731), .Y(n302) );
  INVX1 U9983 ( .A(n302), .Y(n7801) );
  AND2X1 U9984 ( .A(n10097), .B(n10079), .Y(n1477) );
  INVX1 U9985 ( .A(n1477), .Y(n7802) );
  AND2X1 U9986 ( .A(n10592), .B(n10574), .Y(n842) );
  INVX1 U9987 ( .A(n842), .Y(n7803) );
  BUFX2 U9988 ( .A(n11252), .Y(n7804) );
  BUFX2 U9989 ( .A(n11251), .Y(n7805) );
  BUFX2 U9990 ( .A(n1539), .Y(n7806) );
  OR2X1 U9991 ( .A(CircularBuffer_len_write_assig_reg_1634[22]), .B(
        CircularBuffer_len_write_assig_reg_1634[21]), .Y(n1546) );
  INVX1 U9992 ( .A(n1546), .Y(n7807) );
  BUFX2 U9993 ( .A(n817), .Y(n7808) );
  OR2X1 U9994 ( .A(CircularBuffer_len_write_assig_2_reg_1729[22]), .B(
        CircularBuffer_len_write_assig_2_reg_1729[21]), .Y(n824) );
  INVX1 U9995 ( .A(n824), .Y(n7809) );
  AND2X1 U9996 ( .A(n10577), .B(n10578), .Y(n861) );
  INVX1 U9997 ( .A(n861), .Y(n7810) );
  AND2X1 U9998 ( .A(n10604), .B(n10576), .Y(n862) );
  INVX1 U9999 ( .A(n862), .Y(n7811) );
  BUFX2 U10000 ( .A(n860), .Y(n7812) );
  AND2X1 U10001 ( .A(n10489), .B(n10491), .Y(n311) );
  INVX1 U10002 ( .A(n311), .Y(n7813) );
  AND2X1 U10003 ( .A(n10483), .B(n10485), .Y(n312) );
  INVX1 U10004 ( .A(n312), .Y(n7814) );
  BUFX2 U10005 ( .A(n310), .Y(n7815) );
  AND2X1 U10006 ( .A(n9913), .B(n9828), .Y(n2057) );
  INVX1 U10007 ( .A(n2057), .Y(n7816) );
  AND2X1 U10008 ( .A(n9915), .B(n9914), .Y(n2058) );
  INVX1 U10009 ( .A(n2058), .Y(n7817) );
  BUFX2 U10010 ( .A(n2056), .Y(n7818) );
  AND2X1 U10011 ( .A(n10124), .B(n10125), .Y(n3191) );
  INVX1 U10012 ( .A(n3191), .Y(n7819) );
  AND2X1 U10013 ( .A(n10122), .B(n10123), .Y(n3192) );
  INVX1 U10014 ( .A(n3192), .Y(n7820) );
  BUFX2 U10015 ( .A(n3190), .Y(n7821) );
  AND2X1 U10016 ( .A(n10619), .B(n10620), .Y(n3243) );
  INVX1 U10017 ( .A(n3243), .Y(n7822) );
  AND2X1 U10018 ( .A(n10617), .B(n10618), .Y(n3244) );
  INVX1 U10019 ( .A(n3244), .Y(n7823) );
  BUFX2 U10020 ( .A(n3242), .Y(n7824) );
  AND2X1 U10021 ( .A(n373), .B(n9933), .Y(N466) );
  INVX1 U10022 ( .A(N466), .Y(n7825) );
  AND2X1 U10023 ( .A(n11205), .B(n8398), .Y(n11206) );
  INVX1 U10024 ( .A(n11206), .Y(n7826) );
  AND2X1 U10025 ( .A(n11175), .B(n8399), .Y(n11176) );
  INVX1 U10026 ( .A(n11176), .Y(n7827) );
  AND2X1 U10027 ( .A(n11218), .B(n8400), .Y(n11219) );
  INVX1 U10028 ( .A(n11219), .Y(n7828) );
  AND2X1 U10029 ( .A(n11188), .B(n8401), .Y(n11189) );
  INVX1 U10030 ( .A(n11189), .Y(n7829) );
  AND2X1 U10031 ( .A(n11208), .B(n8102), .Y(n11209) );
  INVX1 U10032 ( .A(n11209), .Y(n7830) );
  AND2X1 U10033 ( .A(n11178), .B(n8103), .Y(n11179) );
  INVX1 U10034 ( .A(n11179), .Y(n7831) );
  AND2X1 U10035 ( .A(sum_phi_fu_311_p4[31]), .B(n9765), .Y(n11519) );
  INVX1 U10036 ( .A(n11519), .Y(n7832) );
  AND2X1 U10037 ( .A(sum_1_phi_fu_379_p4[31]), .B(n9646), .Y(n11777) );
  INVX1 U10038 ( .A(n11777), .Y(n7833) );
  BUFX2 U10039 ( .A(n11058), .Y(n7834) );
  AND2X1 U10040 ( .A(recentdatapoints_len_load_op_fu_556_p2[12]), .B(n8972), 
        .Y(n1834) );
  INVX1 U10041 ( .A(n1834), .Y(n7835) );
  AND2X1 U10042 ( .A(recentdatapoints_len_load_op_fu_556_p2[25]), .B(n8972), 
        .Y(n1851) );
  INVX1 U10043 ( .A(n1851), .Y(n7836) );
  AND2X1 U10044 ( .A(recentdatapoints_len_load_op_fu_556_p2[29]), .B(n8972), 
        .Y(n1856) );
  INVX1 U10045 ( .A(n1856), .Y(n7837) );
  AND2X1 U10046 ( .A(n8976), .B(n2022), .Y(n2020) );
  INVX1 U10047 ( .A(n2020), .Y(n7838) );
  OR2X1 U10048 ( .A(n8379), .B(recentdatapoints_len_load_op_fu_556_p2[2]), .Y(
        n2022) );
  AND2X1 U10049 ( .A(n9935), .B(tmp_33_i_fu_786_p2[4]), .Y(n1708) );
  INVX1 U10050 ( .A(n1708), .Y(n7839) );
  AND2X1 U10051 ( .A(n10243), .B(tmp_33_i1_fu_1099_p2[3]), .Y(n1223) );
  INVX1 U10052 ( .A(n1223), .Y(n7840) );
  BUFX2 U10053 ( .A(n2190), .Y(n7841) );
  OR2X1 U10054 ( .A(i_11_fu_1179_p2[3]), .B(n8640), .Y(n8849) );
  AND2X1 U10055 ( .A(ap_CS_fsm[13]), .B(ap_rst_n), .Y(
        \Decision_AXILiteS_s_axi_U/n627 ) );
  INVX1 U10056 ( .A(\Decision_AXILiteS_s_axi_U/n627 ), .Y(n7842) );
  AND2X1 U10057 ( .A(VCaptureThresh_loc_reg_298[15]), .B(n8113), .Y(n12105) );
  INVX1 U10058 ( .A(n12105), .Y(n7843) );
  AND2X1 U10059 ( .A(ACaptureThresh_loc_reg_288[15]), .B(n8114), .Y(n11641) );
  INVX1 U10060 ( .A(n11641), .Y(n7844) );
  AND2X1 U10061 ( .A(VCaptureThresh_loc_reg_298[7]), .B(n8111), .Y(n12125) );
  INVX1 U10062 ( .A(n12125), .Y(n7845) );
  AND2X1 U10063 ( .A(ACaptureThresh_loc_reg_288[7]), .B(n8112), .Y(n11661) );
  INVX1 U10064 ( .A(n11661), .Y(n7846) );
  BUFX2 U10065 ( .A(\Decision_AXILiteS_s_axi_U/n616 ), .Y(n7847) );
  BUFX2 U10066 ( .A(n11410), .Y(n7848) );
  BUFX2 U10067 ( .A(n11408), .Y(n7849) );
  BUFX2 U10068 ( .A(n11407), .Y(n7850) );
  BUFX2 U10069 ( .A(n11315), .Y(n7851) );
  BUFX2 U10070 ( .A(n11316), .Y(n7852) );
  BUFX2 U10071 ( .A(n11263), .Y(n7853) );
  BUFX2 U10072 ( .A(n11264), .Y(n7854) );
  BUFX2 U10073 ( .A(\Decision_AXILiteS_s_axi_U/n570 ), .Y(n7855) );
  AND2X1 U10074 ( .A(recentdatapoints_data_q0[9]), .B(n8868), .Y(n400) );
  INVX1 U10075 ( .A(n400), .Y(n7856) );
  AND2X1 U10076 ( .A(recentdatapoints_data_q0[5]), .B(n8869), .Y(n408) );
  INVX1 U10077 ( .A(n408), .Y(n7857) );
  AND2X1 U10078 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[12]), 
        .Y(n465) );
  INVX1 U10079 ( .A(n465), .Y(n7858) );
  AND2X1 U10080 ( .A(CircularBuffer_len_read_assign_fu_772_p2[10]), .B(n3151), 
        .Y(n2774) );
  INVX1 U10081 ( .A(n2774), .Y(n7859) );
  AND2X1 U10082 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[10]), .B(
        n3149), .Y(n2281) );
  INVX1 U10083 ( .A(n2281), .Y(n7860) );
  AND2X1 U10084 ( .A(CircularBuffer_len_read_assign_fu_772_p2[9]), .B(n3151), 
        .Y(n2776) );
  INVX1 U10085 ( .A(n2776), .Y(n7861) );
  AND2X1 U10086 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[9]), .B(n3149), .Y(n2283) );
  INVX1 U10087 ( .A(n2283), .Y(n7862) );
  AND2X1 U10088 ( .A(CircularBuffer_len_read_assign_fu_772_p2[19]), .B(n8919), 
        .Y(n2756) );
  INVX1 U10089 ( .A(n2756), .Y(n7863) );
  AND2X1 U10090 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[19]), .B(
        n8921), .Y(n2263) );
  INVX1 U10091 ( .A(n2263), .Y(n7864) );
  AND2X1 U10092 ( .A(n8882), .B(\Decision_AXILiteS_s_axi_U/n384 ), .Y(
        \Decision_AXILiteS_s_axi_U/n484 ) );
  INVX1 U10093 ( .A(\Decision_AXILiteS_s_axi_U/n484 ), .Y(n7865) );
  AND2X1 U10094 ( .A(\Decision_AXILiteS_s_axi_U/n397 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n386 ) );
  INVX1 U10095 ( .A(\Decision_AXILiteS_s_axi_U/n386 ), .Y(n7866) );
  BUFX2 U10096 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n40 ), .Y(n7867) );
  BUFX2 U10097 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n42 ), .Y(n7868) );
  BUFX2 U10098 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n38 ), .Y(n7869) );
  AND2X1 U10099 ( .A(\Decision_AXILiteS_s_axi_U/n385 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n419 ) );
  INVX1 U10100 ( .A(\Decision_AXILiteS_s_axi_U/n419 ), .Y(n7870) );
  AND2X1 U10101 ( .A(\Decision_AXILiteS_s_axi_U/n353 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n545 ) );
  INVX1 U10102 ( .A(\Decision_AXILiteS_s_axi_U/n545 ), .Y(n7871) );
  AND2X1 U10103 ( .A(p_tmp_i_reg_1556[3]), .B(n8664), .Y(n8854) );
  OR2X1 U10104 ( .A(CircularBuffer_len_read_assign_1_reg_1616[30]), .B(n8834), 
        .Y(n8853) );
  AND2X1 U10105 ( .A(s_axi_AXILiteS_ARVALID), .B(s_axi_AXILiteS_ARREADY), .Y(
        \Decision_AXILiteS_s_axi_U/n630 ) );
  AND2X1 U10106 ( .A(a_length[1]), .B(n8951), .Y(n3124) );
  INVX1 U10107 ( .A(n3124), .Y(n7872) );
  AND2X1 U10108 ( .A(a_length[13]), .B(n8952), .Y(n3100) );
  INVX1 U10109 ( .A(n3100), .Y(n7873) );
  AND2X1 U10110 ( .A(v_length[7]), .B(n8954), .Y(n2984) );
  INVX1 U10111 ( .A(n2984), .Y(n7874) );
  AND2X1 U10112 ( .A(v_length[23]), .B(n8955), .Y(n2952) );
  INVX1 U10113 ( .A(n2952), .Y(n7875) );
  AND2X1 U10114 ( .A(a_flip[1]), .B(n8953), .Y(n2867) );
  INVX1 U10115 ( .A(n2867), .Y(n7876) );
  AND2X1 U10116 ( .A(p_tmp_i_reg_1556[30]), .B(n8979), .Y(n1922) );
  INVX1 U10117 ( .A(n1922), .Y(n7877) );
  AND2X1 U10118 ( .A(p_tmp_i_reg_1556[18]), .B(n8980), .Y(n1898) );
  INVX1 U10119 ( .A(n1898), .Y(n7878) );
  AND2X1 U10120 ( .A(p_tmp_i_reg_1556[6]), .B(n8977), .Y(n1874) );
  INVX1 U10121 ( .A(n1874), .Y(n7879) );
  AND2X1 U10122 ( .A(recentVBools_head_i[18]), .B(n9010), .Y(n1750) );
  INVX1 U10123 ( .A(n1750), .Y(n7880) );
  AND2X1 U10124 ( .A(recentVBools_head_i[25]), .B(n9009), .Y(n1729) );
  INVX1 U10125 ( .A(n1729), .Y(n7881) );
  AND2X1 U10126 ( .A(ap_CS_fsm[2]), .B(recentVBools_head_i[2]), .Y(n1699) );
  INVX1 U10127 ( .A(n1699), .Y(n7882) );
  AND2X1 U10128 ( .A(n8991), .B(CircularBuffer_len_read_assign_1_fu_778_p3[2]), 
        .Y(n1643) );
  INVX1 U10129 ( .A(n1643), .Y(n7883) );
  BUFX2 U10130 ( .A(n2825), .Y(n7884) );
  BUFX2 U10131 ( .A(n2805), .Y(n7885) );
  AND2X1 U10132 ( .A(CircularBuffer_len_write_assig_fu_817_p2[30]), .B(n1646), 
        .Y(n1558) );
  INVX1 U10133 ( .A(n1558), .Y(n7886) );
  AND2X1 U10134 ( .A(CircularBuffer_sum_read_assign_reg_1610[25]), .B(n9006), 
        .Y(n1416) );
  INVX1 U10135 ( .A(n1416), .Y(n7887) );
  AND2X1 U10136 ( .A(CircularBuffer_sum_read_assign_reg_1610[29]), .B(n9007), 
        .Y(n1408) );
  INVX1 U10137 ( .A(n1408), .Y(n7888) );
  AND2X1 U10138 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[1]), .Y(n2692) );
  INVX1 U10139 ( .A(n2692), .Y(n7889) );
  AND2X1 U10140 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[16]), .Y(n2632) );
  INVX1 U10141 ( .A(n2632), .Y(n7890) );
  BUFX2 U10142 ( .A(n2700), .Y(n7891) );
  AND2X1 U10143 ( .A(n9012), .B(sum_phi_fu_311_p4[31]), .Y(n2571) );
  INVX1 U10144 ( .A(n2571), .Y(n7892) );
  AND2X1 U10145 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[23]), .B(n9031), 
        .Y(n1386) );
  INVX1 U10146 ( .A(n1386), .Y(n7893) );
  AND2X1 U10147 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[18]), .B(n9040), 
        .Y(n1303) );
  INVX1 U10148 ( .A(n1303), .Y(n7894) );
  AND2X1 U10149 ( .A(recentABools_head_i[23]), .B(n9039), .Y(n1288) );
  INVX1 U10150 ( .A(n1288), .Y(n7895) );
  AND2X1 U10151 ( .A(recentABools_head_i[28]), .B(n9038), .Y(n1276) );
  INVX1 U10152 ( .A(n1276), .Y(n7896) );
  AND2X1 U10153 ( .A(recentABools_head_i[1]), .B(ap_CS_fsm[7]), .Y(n1210) );
  INVX1 U10154 ( .A(n1210), .Y(n7897) );
  AND2X1 U10155 ( .A(tmp_5_fu_726_p2[1]), .B(n8992), .Y(n1204) );
  INVX1 U10156 ( .A(n1204), .Y(n7898) );
  AND2X1 U10157 ( .A(VbeatFallDelay[15]), .B(n9036), .Y(n1146) );
  INVX1 U10158 ( .A(n1146), .Y(n7899) );
  AND2X1 U10159 ( .A(tmp_5_fu_726_p2[17]), .B(n8993), .Y(n1140) );
  INVX1 U10160 ( .A(n1140), .Y(n7900) );
  AND2X1 U10161 ( .A(VbeatFallDelay_new_1_reg_342[23]), .B(n9013), .Y(n2180)
         );
  INVX1 U10162 ( .A(n2180), .Y(n7901) );
  AND2X1 U10163 ( .A(VbeatFallDelay[24]), .B(n9035), .Y(n1110) );
  INVX1 U10164 ( .A(n1110), .Y(n7902) );
  AND2X1 U10165 ( .A(VbeatFallDelay_new_1_reg_342[31]), .B(n9013), .Y(n2188)
         );
  INVX1 U10166 ( .A(n2188), .Y(n7903) );
  AND2X1 U10167 ( .A(tmp_4_fu_716_p2[3]), .B(n8994), .Y(n1068) );
  INVX1 U10168 ( .A(n1068), .Y(n7904) );
  AND2X1 U10169 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[6]), .Y(n2560) );
  INVX1 U10170 ( .A(n2560), .Y(n7905) );
  AND2X1 U10171 ( .A(VbeatDelay[8]), .B(n9033), .Y(n1051) );
  INVX1 U10172 ( .A(n1051), .Y(n7906) );
  AND2X1 U10173 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[18]), .Y(n2548) );
  INVX1 U10174 ( .A(n2548), .Y(n7907) );
  AND2X1 U10175 ( .A(tmp_4_fu_716_p2[22]), .B(n8995), .Y(n1006) );
  INVX1 U10176 ( .A(n1006), .Y(n7908) );
  AND2X1 U10177 ( .A(VbeatDelay[24]), .B(n9032), .Y(n997) );
  INVX1 U10178 ( .A(n997), .Y(n7909) );
  AND2X1 U10179 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[27]), .Y(n2539) );
  INVX1 U10180 ( .A(n2539), .Y(n7910) );
  AND2X1 U10181 ( .A(VbeatDelay[29]), .B(n9034), .Y(n979) );
  INVX1 U10182 ( .A(n979), .Y(n7911) );
  BUFX2 U10183 ( .A(n2325), .Y(n7912) );
  AND2X1 U10184 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[20]), .Y(n2486) );
  INVX1 U10185 ( .A(n2486), .Y(n7913) );
  BUFX2 U10186 ( .A(n2313), .Y(n7914) );
  AND2X1 U10187 ( .A(n9017), .B(CircularBuffer_len_read_assign_3_fu_1091_p3[3]), .Y(n966) );
  INVX1 U10188 ( .A(n966), .Y(n7915) );
  AND2X1 U10189 ( .A(n2401), .B(n9019), .Y(n927) );
  INVX1 U10190 ( .A(n927), .Y(n7916) );
  BUFX2 U10191 ( .A(n2394), .Y(n7917) );
  BUFX2 U10192 ( .A(n2372), .Y(n7918) );
  BUFX2 U10193 ( .A(n2346), .Y(n7919) );
  AND2X1 U10194 ( .A(CircularBuffer_len_write_assig_2_fu_1142_p2[30]), .B(n970), .Y(n882) );
  INVX1 U10195 ( .A(n882), .Y(n7920) );
  AND2X1 U10196 ( .A(tmp_3_fu_706_p2[4]), .B(n8996), .Y(n779) );
  INVX1 U10197 ( .A(n779), .Y(n7921) );
  AND2X1 U10198 ( .A(AbeatDelay[5]), .B(n8896), .Y(n773) );
  INVX1 U10199 ( .A(n773), .Y(n7922) );
  AND2X1 U10200 ( .A(AbeatDelay_new_reg_394[6]), .B(n9041), .Y(n2228) );
  INVX1 U10201 ( .A(n2228), .Y(n7923) );
  AND2X1 U10202 ( .A(AbeatDelay_new_reg_394[18]), .B(n9041), .Y(n2216) );
  INVX1 U10203 ( .A(n2216), .Y(n7924) );
  AND2X1 U10204 ( .A(tmp_3_fu_706_p2[28]), .B(n8997), .Y(n698) );
  INVX1 U10205 ( .A(n698), .Y(n7925) );
  AND2X1 U10206 ( .A(AbeatDelay_new_reg_394[29]), .B(n9041), .Y(n2205) );
  INVX1 U10207 ( .A(n2205), .Y(n7926) );
  AND2X1 U10208 ( .A(tmp_3_fu_706_p2[31]), .B(ap_CS_fsm[4]), .Y(n688) );
  INVX1 U10209 ( .A(n688), .Y(n7927) );
  AND2X1 U10210 ( .A(AstimDelay[4]), .B(n8896), .Y(n671) );
  INVX1 U10211 ( .A(n671), .Y(n7928) );
  AND2X1 U10212 ( .A(tmp_6_fu_497_p3[7]), .B(n8967), .Y(n663) );
  INVX1 U10213 ( .A(n663), .Y(n7929) );
  AND2X1 U10214 ( .A(AstimDelay[21]), .B(n8896), .Y(n620) );
  INVX1 U10215 ( .A(n620), .Y(n7930) );
  AND2X1 U10216 ( .A(tmp_6_fu_497_p3[25]), .B(n8966), .Y(n609) );
  INVX1 U10217 ( .A(n609), .Y(n7931) );
  AND2X1 U10218 ( .A(VstimDelay[7]), .B(n10670), .Y(n562) );
  INVX1 U10219 ( .A(n562), .Y(n7932) );
  AND2X1 U10220 ( .A(tmp_7_fu_511_p3[10]), .B(n8965), .Y(n554) );
  INVX1 U10221 ( .A(n554), .Y(n7933) );
  AND2X1 U10222 ( .A(VstimDelay[23]), .B(n10670), .Y(n514) );
  INVX1 U10223 ( .A(n514), .Y(n7934) );
  AND2X1 U10224 ( .A(tmp_7_fu_511_p3[30]), .B(n8964), .Y(n494) );
  INVX1 U10225 ( .A(n494), .Y(n7935) );
  AND2X1 U10226 ( .A(VstimDelay[31]), .B(n8896), .Y(n486) );
  INVX1 U10227 ( .A(n486), .Y(n7936) );
  BUFX2 U10228 ( .A(n2303), .Y(n7937) );
  AND2X1 U10229 ( .A(\Decision_AXILiteS_s_axi_U/n358 ), .B(
        \Decision_AXILiteS_s_axi_U/n351 ), .Y(\Decision_AXILiteS_s_axi_U/n357 ) );
  INVX1 U10230 ( .A(\Decision_AXILiteS_s_axi_U/n357 ), .Y(n7938) );
  AND2X1 U10231 ( .A(\Decision_AXILiteS_s_axi_U/n356 ), .B(n8411), .Y(
        \Decision_AXILiteS_s_axi_U/n461 ) );
  INVX1 U10232 ( .A(\Decision_AXILiteS_s_axi_U/n461 ), .Y(n7939) );
  AND2X1 U10233 ( .A(s_axi_AXILiteS_AWADDR[5]), .B(n8652), .Y(
        \Decision_AXILiteS_s_axi_U/n640 ) );
  INVX1 U10234 ( .A(\Decision_AXILiteS_s_axi_U/n640 ), .Y(n7940) );
  AND2X1 U10235 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[6]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n391 )
         );
  INVX1 U10236 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n391 ), 
        .Y(n7941) );
  AND2X1 U10237 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[3]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n420 )
         );
  INVX1 U10238 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n420 ), 
        .Y(n7942) );
  AND2X1 U10239 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[9]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n432 )
         );
  INVX1 U10240 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n432 ), 
        .Y(n7943) );
  AND2X1 U10241 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[2]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n452 )
         );
  INVX1 U10242 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n452 ), 
        .Y(n7944) );
  AND2X1 U10243 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[8]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n464 )
         );
  INVX1 U10244 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n464 ), 
        .Y(n7945) );
  AND2X1 U10245 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[5]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n492 )
         );
  INVX1 U10246 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n492 ), 
        .Y(n7946) );
  AND2X1 U10247 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[11]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n504 )
         );
  INVX1 U10248 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n504 ), 
        .Y(n7947) );
  AND2X1 U10249 ( .A(n9467), .B(data_read_reg_1495[4]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n524 )
         );
  INVX1 U10250 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n524 ), 
        .Y(n7948) );
  AND2X1 U10251 ( .A(n9467), .B(data_read_reg_1495[10]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n536 )
         );
  INVX1 U10252 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n536 ), 
        .Y(n7949) );
  AND2X1 U10253 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][4] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n559 )
         );
  INVX1 U10254 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n559 ), 
        .Y(n7950) );
  AND2X1 U10255 ( .A(n9468), .B(data_read_reg_1495[13]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n610 )
         );
  INVX1 U10256 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n610 ), 
        .Y(n7951) );
  AND2X1 U10257 ( .A(n9469), .B(data_read_reg_1495[12]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n642 )
         );
  INVX1 U10258 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n642 ), 
        .Y(n7952) );
  AND2X1 U10259 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][7] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n660 )
         );
  INVX1 U10260 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n660 ), 
        .Y(n7953) );
  AND2X1 U10261 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][6] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n678 )
         );
  INVX1 U10262 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n678 ), 
        .Y(n7954) );
  AND2X1 U10263 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][9] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n699 )
         );
  INVX1 U10264 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n699 ), 
        .Y(n7955) );
  AND2X1 U10265 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][8] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n715 )
         );
  INVX1 U10266 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n715 ), 
        .Y(n7956) );
  AND2X1 U10267 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][11] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n735 )
         );
  INVX1 U10268 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n735 ), 
        .Y(n7957) );
  AND2X1 U10269 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][10] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n751 )
         );
  INVX1 U10270 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n751 ), 
        .Y(n7958) );
  AND2X1 U10271 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][1] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n759 )
         );
  INVX1 U10272 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n759 ), 
        .Y(n7959) );
  AND2X1 U10273 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][13] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n771 )
         );
  INVX1 U10274 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n771 ), 
        .Y(n7960) );
  AND2X1 U10275 ( .A(n9466), .B(data_read_reg_1495[15]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n806 )
         );
  INVX1 U10276 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n806 ), 
        .Y(n7961) );
  AND2X1 U10277 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][0] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n809 )
         );
  INVX1 U10278 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n809 ), 
        .Y(n7962) );
  AND2X1 U10279 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][12] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n821 )
         );
  INVX1 U10280 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n821 ), 
        .Y(n7963) );
  AND2X1 U10281 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][15] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n842 )
         );
  INVX1 U10282 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n842 ), 
        .Y(n7964) );
  AND2X1 U10283 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][14] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n858 )
         );
  INVX1 U10284 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n858 ), 
        .Y(n7965) );
  AND2X1 U10285 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[14]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n890 )
         );
  INVX1 U10286 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n890 ), 
        .Y(n7966) );
  AND2X1 U10287 ( .A(
        \recentABools_data_U/Decision_recentVBools_data_ram_U/n141 ), .B(n8405), .Y(\recentABools_data_U/Decision_recentVBools_data_ram_U/n11 ) );
  INVX1 U10288 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n11 ), .Y(n7967) );
  AND2X1 U10289 ( .A(sum_reg_308[8]), .B(n8929), .Y(n2666) );
  INVX1 U10290 ( .A(n2666), .Y(n7968) );
  AND2X1 U10291 ( .A(n429), .B(n397), .Y(n430) );
  INVX1 U10292 ( .A(n430), .Y(n7969) );
  AND2X1 U10293 ( .A(tmp_29_i_fu_752_p2[2]), .B(n8920), .Y(n3162) );
  INVX1 U10294 ( .A(n3162), .Y(n7970) );
  AND2X1 U10295 ( .A(tmp_29_i1_fu_1065_p2[2]), .B(n8922), .Y(n3214) );
  INVX1 U10296 ( .A(n3214), .Y(n7971) );
  AND2X1 U10297 ( .A(tmp_29_i_fu_752_p2[0]), .B(n8920), .Y(n3184) );
  INVX1 U10298 ( .A(n3184), .Y(n7972) );
  AND2X1 U10299 ( .A(tmp_29_i1_fu_1065_p2[0]), .B(n8922), .Y(n3236) );
  INVX1 U10300 ( .A(n3236), .Y(n7973) );
  AND2X1 U10301 ( .A(N505), .B(ap_CS_fsm[12]), .Y(n489) );
  INVX1 U10302 ( .A(n489), .Y(n7974) );
  AND2X1 U10303 ( .A(sum_reg_308[29]), .B(n8929), .Y(n2582) );
  INVX1 U10304 ( .A(n2582), .Y(n7975) );
  AND2X1 U10305 ( .A(sum_1_reg_376[29]), .B(n8930), .Y(n2524) );
  INVX1 U10306 ( .A(n2524), .Y(n7976) );
  AND2X1 U10307 ( .A(sum_reg_308[18]), .B(n8929), .Y(n2626) );
  INVX1 U10308 ( .A(n2626), .Y(n7977) );
  AND2X1 U10309 ( .A(sum_1_reg_376[22]), .B(n8930), .Y(n2496) );
  INVX1 U10310 ( .A(n2496), .Y(n7978) );
  INVX1 U10311 ( .A(n3854), .Y(n7979) );
  AND2X1 U10312 ( .A(CircularBuffer_head_i_read_ass_reg_1624[1]), .B(n9008), 
        .Y(n1696) );
  INVX1 U10313 ( .A(n1696), .Y(n7980) );
  INVX1 U10314 ( .A(n3650), .Y(n7981) );
  AND2X1 U10315 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[1]), .B(n9037), 
        .Y(n1213) );
  INVX1 U10316 ( .A(n1213), .Y(n7982) );
  INVX1 U10317 ( .A(n4622), .Y(n7983) );
  AND2X1 U10318 ( .A(ACaptureThresh_loc_reg_288[12]), .B(n8970), .Y(n3038) );
  INVX1 U10319 ( .A(n3038), .Y(n7984) );
  BUFX2 U10320 ( .A(n3037), .Y(n7985) );
  INVX1 U10321 ( .A(n4609), .Y(n7986) );
  AND2X1 U10322 ( .A(ACaptureThresh_loc_reg_288[25]), .B(n8971), .Y(n3012) );
  INVX1 U10323 ( .A(n3012), .Y(n7987) );
  BUFX2 U10324 ( .A(n3011), .Y(n7988) );
  INVX1 U10325 ( .A(n4564), .Y(n7989) );
  AND2X1 U10326 ( .A(VCaptureThresh_loc_reg_298[6]), .B(n8970), .Y(n2922) );
  INVX1 U10327 ( .A(n2922), .Y(n7990) );
  BUFX2 U10328 ( .A(n2921), .Y(n7991) );
  INVX1 U10329 ( .A(n4551), .Y(n7992) );
  AND2X1 U10330 ( .A(VCaptureThresh_loc_reg_298[19]), .B(n8969), .Y(n2896) );
  INVX1 U10331 ( .A(n2896), .Y(n7993) );
  BUFX2 U10332 ( .A(n2895), .Y(n7994) );
  INVX1 U10333 ( .A(n4539), .Y(n7995) );
  AND2X1 U10334 ( .A(VCaptureThresh_loc_reg_298[31]), .B(n8968), .Y(n2871) );
  INVX1 U10335 ( .A(n2871), .Y(n7996) );
  BUFX2 U10336 ( .A(n2870), .Y(n7997) );
  OR2X1 U10337 ( .A(VbeatFallDelay_new_1_reg_342[20]), .B(
        VbeatFallDelay_new_1_reg_342[19]), .Y(n11905) );
  INVX1 U10338 ( .A(n11905), .Y(n7998) );
  OR2X1 U10339 ( .A(n9320), .B(n8383), .Y(\Decision_AXILiteS_s_axi_U/n334 ) );
  INVX1 U10340 ( .A(\Decision_AXILiteS_s_axi_U/n334 ), .Y(n7999) );
  AND2X1 U10341 ( .A(tmp_6_reg_1538[29]), .B(n9638), .Y(n11977) );
  INVX1 U10342 ( .A(n11977), .Y(n8000) );
  AND2X1 U10343 ( .A(tmp_7_reg_1544[29]), .B(n9755), .Y(n12066) );
  INVX1 U10344 ( .A(n12066), .Y(n8001) );
  AND2X1 U10345 ( .A(VbeatDelay_new_1_reg_326[13]), .B(n10705), .Y(n11098) );
  INVX1 U10346 ( .A(n11098), .Y(n8002) );
  AND2X1 U10347 ( .A(VbeatDelay_new_1_reg_326[29]), .B(n10443), .Y(n11869) );
  INVX1 U10348 ( .A(n11869), .Y(n8003) );
  BUFX2 U10349 ( .A(n11909), .Y(n8004) );
  BUFX2 U10350 ( .A(n11910), .Y(n8005) );
  OR2X1 U10351 ( .A(CircularBuffer_head_i_read_ass_reg_1624[7]), .B(n11310), 
        .Y(n11312) );
  INVX1 U10352 ( .A(n11312), .Y(n8006) );
  AND2X1 U10353 ( .A(CircularBuffer_head_i_read_ass_reg_1624[7]), .B(n11310), 
        .Y(n11311) );
  INVX1 U10354 ( .A(n11311), .Y(n8007) );
  OR2X1 U10355 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[7]), .B(n11258), 
        .Y(n11260) );
  INVX1 U10356 ( .A(n11260), .Y(n8008) );
  AND2X1 U10357 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[7]), .B(n11258), 
        .Y(n11259) );
  INVX1 U10358 ( .A(n11259), .Y(n8009) );
  BUFX2 U10359 ( .A(n12032), .Y(n8010) );
  BUFX2 U10360 ( .A(n12029), .Y(n8011) );
  BUFX2 U10361 ( .A(n11111), .Y(n8012) );
  BUFX2 U10362 ( .A(n11108), .Y(n8013) );
  OR2X1 U10363 ( .A(VbeatDelay_new_1_reg_326[11]), .B(
        VbeatDelay_new_1_reg_326[10]), .Y(n318) );
  INVX1 U10364 ( .A(n318), .Y(n8014) );
  OR2X1 U10365 ( .A(recentdatapoints_len[9]), .B(recentdatapoints_len[8]), .Y(
        n2045) );
  INVX1 U10366 ( .A(n2045), .Y(n8015) );
  OR2X1 U10367 ( .A(recentdatapoints_len[10]), .B(recentdatapoints_len[0]), 
        .Y(n2036) );
  INVX1 U10368 ( .A(n2036), .Y(n8016) );
  OR2X1 U10369 ( .A(p_tmp_i_fu_587_p3[9]), .B(p_tmp_i_fu_587_p3[8]), .Y(n1949)
         );
  INVX1 U10370 ( .A(n1949), .Y(n8017) );
  OR2X1 U10371 ( .A(VbeatDelay_new_1_reg_326[4]), .B(
        VbeatDelay_new_1_reg_326[3]), .Y(n338) );
  INVX1 U10372 ( .A(n338), .Y(n8018) );
  AND2X1 U10373 ( .A(n10575), .B(n10603), .Y(n870) );
  INVX1 U10374 ( .A(n870), .Y(n8019) );
  AND2X1 U10375 ( .A(vflip[5]), .B(vflip[4]), .Y(n436) );
  INVX1 U10376 ( .A(n436), .Y(n8020) );
  AND2X1 U10377 ( .A(aflip[5]), .B(aflip[4]), .Y(n478) );
  INVX1 U10378 ( .A(n478), .Y(n8021) );
  AND2X1 U10379 ( .A(n10517), .B(n10521), .Y(n342) );
  INVX1 U10380 ( .A(n342), .Y(n8022) );
  AND2X1 U10381 ( .A(n10082), .B(n10083), .Y(n1496) );
  INVX1 U10382 ( .A(n1496), .Y(n8023) );
  AND2X1 U10383 ( .A(n10109), .B(n10081), .Y(n1497) );
  INVX1 U10384 ( .A(n1497), .Y(n8024) );
  BUFX2 U10385 ( .A(n1495), .Y(n8025) );
  AND2X1 U10386 ( .A(n9877), .B(n9876), .Y(n1938) );
  INVX1 U10387 ( .A(n1938), .Y(n8026) );
  AND2X1 U10388 ( .A(n9879), .B(n9878), .Y(n1939) );
  INVX1 U10389 ( .A(n1939), .Y(n8027) );
  BUFX2 U10390 ( .A(n1937), .Y(n8028) );
  AND2X1 U10391 ( .A(n9928), .B(n9927), .Y(n2066) );
  INVX1 U10392 ( .A(n2066), .Y(n8029) );
  AND2X1 U10393 ( .A(n9901), .B(n9929), .Y(n2067) );
  INVX1 U10394 ( .A(n2067), .Y(n8030) );
  BUFX2 U10395 ( .A(n2065), .Y(n8031) );
  AND2X1 U10396 ( .A(n10172), .B(n10114), .Y(n3200) );
  INVX1 U10397 ( .A(n3200), .Y(n8032) );
  AND2X1 U10398 ( .A(n10138), .B(n10078), .Y(n3201) );
  INVX1 U10399 ( .A(n3201), .Y(n8033) );
  BUFX2 U10400 ( .A(n3199), .Y(n8034) );
  AND2X1 U10401 ( .A(n10669), .B(n10609), .Y(n3252) );
  INVX1 U10402 ( .A(n3252), .Y(n8035) );
  AND2X1 U10403 ( .A(n10633), .B(n10573), .Y(n3253) );
  INVX1 U10404 ( .A(n3253), .Y(n8036) );
  BUFX2 U10405 ( .A(n3251), .Y(n8037) );
  AND2X1 U10406 ( .A(n10095), .B(n10096), .Y(n1478) );
  INVX1 U10407 ( .A(n1478), .Y(n8038) );
  AND2X1 U10408 ( .A(n10590), .B(n10591), .Y(n843) );
  INVX1 U10409 ( .A(n843), .Y(n8039) );
  AND2X1 U10410 ( .A(n9916), .B(n9915), .Y(n1656) );
  INVX1 U10411 ( .A(n1656), .Y(n8040) );
  AND2X1 U10412 ( .A(n9918), .B(n9917), .Y(n1657) );
  INVX1 U10413 ( .A(n1657), .Y(n8041) );
  BUFX2 U10414 ( .A(n1655), .Y(n8042) );
  BUFX2 U10415 ( .A(n1522), .Y(n8043) );
  OR2X1 U10416 ( .A(CircularBuffer_len_write_assig_reg_1634[26]), .B(
        CircularBuffer_len_write_assig_reg_1634[25]), .Y(n1525) );
  INVX1 U10417 ( .A(n1525), .Y(n8044) );
  BUFX2 U10418 ( .A(n800), .Y(n8045) );
  OR2X1 U10419 ( .A(CircularBuffer_len_write_assig_2_reg_1729[26]), .B(
        CircularBuffer_len_write_assig_2_reg_1729[25]), .Y(n803) );
  INVX1 U10420 ( .A(n803), .Y(n8046) );
  BUFX2 U10421 ( .A(n11250), .Y(n8047) );
  OR2X1 U10422 ( .A(p_tmp_i_reg_1556[11]), .B(p_tmp_i_reg_1556[10]), .Y(n11249) );
  INVX1 U10423 ( .A(n11249), .Y(n8048) );
  AND2X1 U10424 ( .A(n387), .B(n9013), .Y(N461) );
  INVX1 U10425 ( .A(N461), .Y(n8049) );
  AND2X1 U10426 ( .A(n11232), .B(n8406), .Y(n11233) );
  INVX1 U10427 ( .A(n11233), .Y(n8050) );
  AND2X1 U10428 ( .A(n11202), .B(n8407), .Y(n11203) );
  INVX1 U10429 ( .A(n11203), .Y(n8051) );
  AND2X1 U10430 ( .A(n11225), .B(n10072), .Y(n11228) );
  INVX1 U10431 ( .A(n11228), .Y(n8052) );
  AND2X1 U10432 ( .A(n11195), .B(n10537), .Y(n11198) );
  INVX1 U10433 ( .A(n11198), .Y(n8053) );
  AND2X1 U10434 ( .A(n10074), .B(n8391), .Y(n11214) );
  INVX1 U10435 ( .A(n11214), .Y(n8054) );
  AND2X1 U10436 ( .A(n10539), .B(n8392), .Y(n11184) );
  INVX1 U10437 ( .A(n11184), .Y(n8055) );
  AND2X1 U10438 ( .A(n11235), .B(n9898), .Y(n11246) );
  INVX1 U10439 ( .A(n11246), .Y(n8056) );
  AND2X1 U10440 ( .A(recentdatapoints_len_load_op_fu_556_p2[13]), .B(n8972), 
        .Y(n1835) );
  INVX1 U10441 ( .A(n1835), .Y(n8057) );
  AND2X1 U10442 ( .A(recentdatapoints_len_load_op_fu_556_p2[26]), .B(n8972), 
        .Y(n1853) );
  INVX1 U10443 ( .A(n1853), .Y(n8058) );
  AND2X1 U10444 ( .A(recentdatapoints_len_load_op_fu_556_p2[30]), .B(n8972), 
        .Y(n1857) );
  INVX1 U10445 ( .A(n1857), .Y(n8059) );
  AND2X1 U10446 ( .A(n8975), .B(n2017), .Y(n1824) );
  INVX1 U10447 ( .A(n1824), .Y(n8060) );
  OR2X1 U10448 ( .A(n8379), .B(recentdatapoints_len_load_op_fu_556_p2[4]), .Y(
        n2017) );
  AND2X1 U10449 ( .A(n9935), .B(tmp_33_i_fu_786_p2[2]), .Y(n1701) );
  INVX1 U10450 ( .A(n1701), .Y(n8061) );
  AND2X1 U10451 ( .A(n10243), .B(tmp_33_i1_fu_1099_p2[2]), .Y(n1218) );
  INVX1 U10452 ( .A(n1218), .Y(n8062) );
  BUFX2 U10453 ( .A(n11482), .Y(n8063) );
  BUFX2 U10454 ( .A(n11937), .Y(n8064) );
  BUFX2 U10455 ( .A(n12026), .Y(n8065) );
  BUFX2 U10456 ( .A(n11829), .Y(n8066) );
  BUFX2 U10457 ( .A(n11740), .Y(n8067) );
  BUFX2 U10458 ( .A(n12235), .Y(n8068) );
  AND2X1 U10459 ( .A(n364), .B(n9933), .Y(n367) );
  INVX1 U10460 ( .A(n367), .Y(n8069) );
  AND2X1 U10461 ( .A(a_thresh[15]), .B(n9479), .Y(n11590) );
  INVX1 U10462 ( .A(n11590), .Y(n8070) );
  AND2X1 U10463 ( .A(tmp_6_reg_1538[31]), .B(n9646), .Y(n11974) );
  INVX1 U10464 ( .A(n11974), .Y(n8071) );
  AND2X1 U10465 ( .A(tmp_7_reg_1544[31]), .B(n9765), .Y(n12063) );
  INVX1 U10466 ( .A(n12063), .Y(n8072) );
  AND2X1 U10467 ( .A(AbeatDelay_new_reg_394[27]), .B(n10523), .Y(n11135) );
  INVX1 U10468 ( .A(n11135), .Y(n8073) );
  AND2X1 U10469 ( .A(AbeatDelay_new_reg_394[15]), .B(n10491), .Y(n11095) );
  INVX1 U10470 ( .A(n11095), .Y(n8074) );
  AND2X1 U10471 ( .A(AbeatDelay_new_reg_394[11]), .B(n10480), .Y(n11089) );
  INVX1 U10472 ( .A(n11089), .Y(n8075) );
  AND2X1 U10473 ( .A(VbeatDelay_new_1_reg_326[31]), .B(n10449), .Y(n11866) );
  INVX1 U10474 ( .A(n11866), .Y(n8076) );
  AND2X1 U10475 ( .A(VCaptureThresh_loc_reg_298[11]), .B(n8398), .Y(n12099) );
  INVX1 U10476 ( .A(n12099), .Y(n8077) );
  AND2X1 U10477 ( .A(ACaptureThresh_loc_reg_288[11]), .B(n8399), .Y(n11635) );
  INVX1 U10478 ( .A(n11635), .Y(n8078) );
  AND2X1 U10479 ( .A(AbeatDelay_new_reg_394[23]), .B(n10512), .Y(n11159) );
  INVX1 U10480 ( .A(n11159), .Y(n8079) );
  AND2X1 U10481 ( .A(AbeatDelay_new_reg_394[19]), .B(n10501), .Y(n11152) );
  INVX1 U10482 ( .A(n11152), .Y(n8080) );
  AND2X1 U10483 ( .A(ACaptureThresh_loc_reg_288[3]), .B(n10746), .Y(n11944) );
  INVX1 U10484 ( .A(n11944), .Y(n8081) );
  AND2X1 U10485 ( .A(VCaptureThresh_loc_reg_298[3]), .B(n10780), .Y(n12033) );
  INVX1 U10486 ( .A(n12033), .Y(n8082) );
  AND2X1 U10487 ( .A(AbeatDelay_new_reg_394[3]), .B(n10459), .Y(n11112) );
  INVX1 U10488 ( .A(n11112), .Y(n8083) );
  AND2X1 U10489 ( .A(AbeatDelay_new_reg_394[7]), .B(n10468), .Y(n11115) );
  INVX1 U10490 ( .A(n11115), .Y(n8084) );
  AND2X1 U10491 ( .A(VCaptureThresh_loc_reg_298[23]), .B(n8400), .Y(n12169) );
  INVX1 U10492 ( .A(n12169), .Y(n8085) );
  AND2X1 U10493 ( .A(ACaptureThresh_loc_reg_288[23]), .B(n8401), .Y(n11705) );
  INVX1 U10494 ( .A(n11705), .Y(n8086) );
  OR2X1 U10495 ( .A(n9540), .B(v_thresh[31]), .Y(n12248) );
  INVX1 U10496 ( .A(n12248), .Y(n8087) );
  OR2X1 U10497 ( .A(n9490), .B(a_thresh[31]), .Y(n11615) );
  INVX1 U10498 ( .A(n11615), .Y(n8088) );
  OR2X1 U10499 ( .A(n10697), .B(VbeatDelay_new_1_reg_326[9]), .Y(n11106) );
  INVX1 U10500 ( .A(n11106), .Y(n8089) );
  BUFX2 U10501 ( .A(n11361), .Y(n8090) );
  BUFX2 U10502 ( .A(n11351), .Y(n8091) );
  BUFX2 U10503 ( .A(n11352), .Y(n8092) );
  BUFX2 U10504 ( .A(n11455), .Y(n8093) );
  BUFX2 U10505 ( .A(n11456), .Y(n8094) );
  BUFX2 U10506 ( .A(n11413), .Y(n8095) );
  BUFX2 U10507 ( .A(n11306), .Y(n8096) );
  BUFX2 U10508 ( .A(n11304), .Y(n8097) );
  BUFX2 U10509 ( .A(n11303), .Y(n8098) );
  BUFX2 U10510 ( .A(n11151), .Y(n8099) );
  BUFX2 U10511 ( .A(n2198), .Y(n8100) );
  AND2X1 U10512 ( .A(recentdatapoints_data_q0[4]), .B(n8869), .Y(n410) );
  INVX1 U10513 ( .A(n410), .Y(n8101) );
  AND2X1 U10514 ( .A(CircularBuffer_len_read_assign_fu_772_p2[14]), .B(n3151), 
        .Y(n2766) );
  INVX1 U10515 ( .A(n2766), .Y(n8102) );
  AND2X1 U10516 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[14]), .B(
        n3149), .Y(n2273) );
  INVX1 U10517 ( .A(n2273), .Y(n8103) );
  OR2X1 U10518 ( .A(n9042), .B(s_axi_AXILiteS_WSTRB[0]), .Y(
        \Decision_AXILiteS_s_axi_U/n565 ) );
  INVX1 U10519 ( .A(\Decision_AXILiteS_s_axi_U/n565 ), .Y(n8104) );
  INVX1 U10520 ( .A(\Decision_AXILiteS_s_axi_U/n607 ), .Y(n8105) );
  BUFX2 U10521 ( .A(\Decision_AXILiteS_s_axi_U/n610 ), .Y(n8106) );
  AND2X1 U10522 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[0]), 
        .Y(n471) );
  INVX1 U10523 ( .A(n471), .Y(n8107) );
  INVX1 U10524 ( .A(recentVBools_data_address0[3]), .Y(n8108) );
  BUFX2 U10525 ( .A(n374), .Y(n8109) );
  BUFX2 U10526 ( .A(n375), .Y(n8110) );
  AND2X1 U10527 ( .A(CircularBuffer_len_read_assign_fu_772_p2[7]), .B(n3151), 
        .Y(n2780) );
  INVX1 U10528 ( .A(n2780), .Y(n8111) );
  AND2X1 U10529 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[7]), .B(n3149), .Y(n2287) );
  INVX1 U10530 ( .A(n2287), .Y(n8112) );
  AND2X1 U10531 ( .A(CircularBuffer_len_read_assign_fu_772_p2[15]), .B(n8919), 
        .Y(n2764) );
  INVX1 U10532 ( .A(n2764), .Y(n8113) );
  AND2X1 U10533 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[15]), .B(
        n8921), .Y(n2271) );
  INVX1 U10534 ( .A(n2271), .Y(n8114) );
  AND2X1 U10535 ( .A(recentdatapoints_data_q0[15]), .B(n8868), .Y(n398) );
  INVX1 U10536 ( .A(n398), .Y(n8115) );
  AND2X1 U10537 ( .A(\Decision_AXILiteS_s_axi_U/n429 ), .B(
        \Decision_AXILiteS_s_axi_U/n384 ), .Y(\Decision_AXILiteS_s_axi_U/n421 ) );
  INVX1 U10538 ( .A(\Decision_AXILiteS_s_axi_U/n421 ), .Y(n8116) );
  BUFX2 U10539 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n38 ), .Y(n8117) );
  BUFX2 U10540 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n44 ), .Y(n8118) );
  BUFX2 U10541 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n40 ), .Y(n8119) );
  AND2X1 U10542 ( .A(\Decision_AXILiteS_s_axi_U/n353 ), .B(n8881), .Y(
        \Decision_AXILiteS_s_axi_U/n398 ) );
  INVX1 U10543 ( .A(\Decision_AXILiteS_s_axi_U/n398 ), .Y(n8120) );
  AND2X1 U10544 ( .A(\Decision_AXILiteS_s_axi_U/n385 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n482 ) );
  INVX1 U10545 ( .A(\Decision_AXILiteS_s_axi_U/n482 ), .Y(n8121) );
  AND2X1 U10546 ( .A(\Decision_AXILiteS_s_axi_U/n397 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n535 ) );
  INVX1 U10547 ( .A(\Decision_AXILiteS_s_axi_U/n535 ), .Y(n8122) );
  OR2X1 U10548 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[30] ), .B(
        n8631), .Y(n8846) );
  AND2X1 U10549 ( .A(a_length[14]), .B(n8952), .Y(n3098) );
  INVX1 U10550 ( .A(n3098), .Y(n8123) );
  AND2X1 U10551 ( .A(v_length[8]), .B(n8954), .Y(n2982) );
  INVX1 U10552 ( .A(n2982), .Y(n8124) );
  AND2X1 U10553 ( .A(v_length[24]), .B(n8955), .Y(n2950) );
  INVX1 U10554 ( .A(n2950), .Y(n8125) );
  AND2X1 U10555 ( .A(a_flip[2]), .B(n8953), .Y(n2865) );
  INVX1 U10556 ( .A(n2865), .Y(n8126) );
  AND2X1 U10557 ( .A(p_tmp_i_reg_1556[26]), .B(n8979), .Y(n1914) );
  INVX1 U10558 ( .A(n1914), .Y(n8127) );
  AND2X1 U10559 ( .A(p_tmp_i_reg_1556[12]), .B(n8980), .Y(n1886) );
  INVX1 U10560 ( .A(n1886), .Y(n8128) );
  AND2X1 U10561 ( .A(p_tmp_i_reg_1556[5]), .B(n8977), .Y(n1872) );
  INVX1 U10562 ( .A(n1872), .Y(n8129) );
  AND2X1 U10563 ( .A(recentVBools_head_i[8]), .B(n9011), .Y(n1780) );
  INVX1 U10564 ( .A(n1780), .Y(n8130) );
  AND2X1 U10565 ( .A(CircularBuffer_head_i_read_ass_reg_1624[19]), .B(n9010), 
        .Y(n1748) );
  INVX1 U10566 ( .A(n1748), .Y(n8131) );
  AND2X1 U10567 ( .A(recentVBools_head_i[26]), .B(n9009), .Y(n1726) );
  INVX1 U10568 ( .A(n1726), .Y(n8132) );
  AND2X1 U10569 ( .A(ap_CS_fsm[2]), .B(recentVBools_head_i[1]), .Y(n1693) );
  INVX1 U10570 ( .A(n1693), .Y(n8133) );
  AND2X1 U10571 ( .A(n2734), .B(n8991), .Y(n1604) );
  INVX1 U10572 ( .A(n1604), .Y(n8134) );
  BUFX2 U10573 ( .A(n2849), .Y(n8135) );
  BUFX2 U10574 ( .A(n2813), .Y(n8136) );
  BUFX2 U10575 ( .A(n2803), .Y(n8137) );
  AND2X1 U10576 ( .A(\recentVBools_data_load_reg_1584[0] ), .B(n9934), .Y(
        n1512) );
  INVX1 U10577 ( .A(n1512), .Y(n8138) );
  AND2X1 U10578 ( .A(CircularBuffer_sum_read_assign_reg_1610[0]), .B(n9008), 
        .Y(n1466) );
  INVX1 U10579 ( .A(n1466), .Y(n8139) );
  AND2X1 U10580 ( .A(CircularBuffer_sum_read_assign_reg_1610[26]), .B(n9006), 
        .Y(n1414) );
  INVX1 U10581 ( .A(n1414), .Y(n8140) );
  AND2X1 U10582 ( .A(CircularBuffer_sum_read_assign_reg_1610[30]), .B(n9007), 
        .Y(n1406) );
  INVX1 U10583 ( .A(n1406), .Y(n8141) );
  AND2X1 U10584 ( .A(n9012), .B(sum_phi_fu_311_p4[0]), .Y(n2696) );
  INVX1 U10585 ( .A(n2696), .Y(n8142) );
  AND2X1 U10586 ( .A(n9012), .B(sum_phi_fu_311_p4[26]), .Y(n2592) );
  INVX1 U10587 ( .A(n2592), .Y(n8143) );
  AND2X1 U10588 ( .A(ap_CS_fsm[7]), .B(sum_phi_fu_311_p4[29]), .Y(n2580) );
  INVX1 U10589 ( .A(n2580), .Y(n8144) );
  AND2X1 U10590 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[13]), .B(n9040), 
        .Y(n1313) );
  INVX1 U10591 ( .A(n1313), .Y(n8145) );
  AND2X1 U10592 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[24]), .B(n9039), 
        .Y(n1287) );
  INVX1 U10593 ( .A(n1287), .Y(n8146) );
  AND2X1 U10594 ( .A(recentABools_head_i[29]), .B(n9038), .Y(n1274) );
  INVX1 U10595 ( .A(n1274), .Y(n8147) );
  AND2X1 U10596 ( .A(VbeatFallDelay[4]), .B(n9037), .Y(n1190) );
  INVX1 U10597 ( .A(n1190), .Y(n8148) );
  AND2X1 U10598 ( .A(tmp_5_fu_726_p2[5]), .B(n8992), .Y(n1188) );
  INVX1 U10599 ( .A(n1188), .Y(n8149) );
  AND2X1 U10600 ( .A(VbeatFallDelay_new_1_reg_342[14]), .B(n9013), .Y(n2171)
         );
  INVX1 U10601 ( .A(n2171), .Y(n8150) );
  AND2X1 U10602 ( .A(VbeatFallDelay[14]), .B(n9036), .Y(n1150) );
  INVX1 U10603 ( .A(n1150), .Y(n8151) );
  AND2X1 U10604 ( .A(VbeatFallDelay_new_1_reg_342[28]), .B(n9013), .Y(n2185)
         );
  INVX1 U10605 ( .A(n2185), .Y(n8152) );
  AND2X1 U10606 ( .A(tmp_4_fu_716_p2[4]), .B(n8994), .Y(n1066) );
  INVX1 U10607 ( .A(n1066), .Y(n8153) );
  AND2X1 U10608 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[7]), .Y(n2559) );
  INVX1 U10609 ( .A(n2559), .Y(n8154) );
  AND2X1 U10610 ( .A(VbeatDelay[13]), .B(n9032), .Y(n1034) );
  INVX1 U10611 ( .A(n1034), .Y(n8155) );
  AND2X1 U10612 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[19]), .Y(n2547) );
  INVX1 U10613 ( .A(n2547), .Y(n8156) );
  AND2X1 U10614 ( .A(tmp_4_fu_716_p2[23]), .B(n8995), .Y(n1003) );
  INVX1 U10615 ( .A(n1003), .Y(n8157) );
  AND2X1 U10616 ( .A(VbeatDelay[25]), .B(n9033), .Y(n993) );
  INVX1 U10617 ( .A(n993), .Y(n8158) );
  AND2X1 U10618 ( .A(n2535), .B(VbeatDelay_new_1_reg_326[30]), .Y(n2536) );
  INVX1 U10619 ( .A(n2536), .Y(n8159) );
  AND2X1 U10620 ( .A(VbeatDelay[30]), .B(n9034), .Y(n976) );
  INVX1 U10621 ( .A(n976), .Y(n8160) );
  AND2X1 U10622 ( .A(VbeatDelay[31]), .B(n9035), .Y(n973) );
  INVX1 U10623 ( .A(n973), .Y(n8161) );
  AND2X1 U10624 ( .A(ap_CS_fsm[12]), .B(sum_1_phi_fu_379_p4[21]), .Y(n2490) );
  INVX1 U10625 ( .A(n2490), .Y(n8162) );
  AND2X1 U10626 ( .A(n9017), .B(CircularBuffer_len_read_assign_3_fu_1091_p3[4]), .Y(n965) );
  INVX1 U10627 ( .A(n965), .Y(n8163) );
  BUFX2 U10628 ( .A(n2352), .Y(n8164) );
  AND2X1 U10629 ( .A(\recentABools_data_load_reg_1700[0] ), .B(n10242), .Y(
        n877) );
  INVX1 U10630 ( .A(n877), .Y(n8165) );
  BUFX2 U10631 ( .A(n2336), .Y(n8166) );
  AND2X1 U10632 ( .A(tmp_3_fu_706_p2[2]), .B(n8993), .Y(n786) );
  INVX1 U10633 ( .A(n786), .Y(n8167) );
  AND2X1 U10634 ( .A(AbeatDelay[6]), .B(n10670), .Y(n770) );
  INVX1 U10635 ( .A(n770), .Y(n8168) );
  AND2X1 U10636 ( .A(AbeatDelay_new_reg_394[9]), .B(n9041), .Y(n2225) );
  INVX1 U10637 ( .A(n2225), .Y(n8169) );
  AND2X1 U10638 ( .A(AbeatDelay[24]), .B(n8896), .Y(n710) );
  INVX1 U10639 ( .A(n710), .Y(n8170) );
  AND2X1 U10640 ( .A(tmp_3_fu_706_p2[29]), .B(n8997), .Y(n694) );
  INVX1 U10641 ( .A(n694), .Y(n8171) );
  AND2X1 U10642 ( .A(AbeatDelay_new_reg_394[30]), .B(n9041), .Y(n2203) );
  INVX1 U10643 ( .A(n2203), .Y(n8172) );
  AND2X1 U10644 ( .A(AbeatDelay_new_reg_394[31]), .B(n9041), .Y(n3146) );
  INVX1 U10645 ( .A(n3146), .Y(n8173) );
  AND2X1 U10646 ( .A(AstimDelay[5]), .B(n8896), .Y(n668) );
  INVX1 U10647 ( .A(n668), .Y(n8174) );
  AND2X1 U10648 ( .A(tmp_6_fu_497_p3[8]), .B(n8967), .Y(n660) );
  INVX1 U10649 ( .A(n660), .Y(n8175) );
  AND2X1 U10650 ( .A(AstimDelay[22]), .B(n8896), .Y(n617) );
  INVX1 U10651 ( .A(n617), .Y(n8176) );
  AND2X1 U10652 ( .A(tmp_6_fu_497_p3[26]), .B(n8966), .Y(n606) );
  INVX1 U10653 ( .A(n606), .Y(n8177) );
  AND2X1 U10654 ( .A(VstimDelay[8]), .B(n8896), .Y(n559) );
  INVX1 U10655 ( .A(n559), .Y(n8178) );
  AND2X1 U10656 ( .A(VstimDelay[22]), .B(n8896), .Y(n517) );
  INVX1 U10657 ( .A(n517), .Y(n8179) );
  AND2X1 U10658 ( .A(tmp_7_fu_511_p3[29]), .B(n8964), .Y(n497) );
  INVX1 U10659 ( .A(n497), .Y(n8180) );
  AND2X1 U10660 ( .A(VstimDelay[30]), .B(n10670), .Y(n493) );
  INVX1 U10661 ( .A(n493), .Y(n8181) );
  AND2X1 U10662 ( .A(s_axi_AXILiteS_AWADDR[6]), .B(n8652), .Y(
        \Decision_AXILiteS_s_axi_U/n641 ) );
  INVX1 U10663 ( .A(\Decision_AXILiteS_s_axi_U/n641 ), .Y(n8182) );
  AND2X1 U10664 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 ), 
        .B(data_read_reg_1495[7]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n393 )
         );
  INVX1 U10665 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n393 ), 
        .Y(n8183) );
  AND2X1 U10666 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[2]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n418 )
         );
  INVX1 U10667 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n418 ), 
        .Y(n8184) );
  AND2X1 U10668 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 ), 
        .B(data_read_reg_1495[8]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n430 )
         );
  INVX1 U10669 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n430 ), 
        .Y(n8185) );
  AND2X1 U10670 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[3]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n454 )
         );
  INVX1 U10671 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n454 ), 
        .Y(n8186) );
  AND2X1 U10672 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 ), 
        .B(data_read_reg_1495[9]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n466 )
         );
  INVX1 U10673 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n466 ), 
        .Y(n8187) );
  AND2X1 U10674 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[4]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n490 )
         );
  INVX1 U10675 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n490 ), 
        .Y(n8188) );
  AND2X1 U10676 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 ), 
        .B(data_read_reg_1495[10]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n502 )
         );
  INVX1 U10677 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n502 ), 
        .Y(n8189) );
  AND2X1 U10678 ( .A(n9467), .B(data_read_reg_1495[5]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n526 )
         );
  INVX1 U10679 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n526 ), 
        .Y(n8190) );
  AND2X1 U10680 ( .A(n9467), .B(data_read_reg_1495[11]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n538 )
         );
  INVX1 U10681 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n538 ), 
        .Y(n8191) );
  AND2X1 U10682 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[5][5] ), .B(n8899), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n561 )
         );
  INVX1 U10683 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n561 ), 
        .Y(n8192) );
  AND2X1 U10684 ( .A(n9468), .B(data_read_reg_1495[12]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n608 )
         );
  INVX1 U10685 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n608 ), 
        .Y(n8193) );
  AND2X1 U10686 ( .A(n9469), .B(data_read_reg_1495[13]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n644 )
         );
  INVX1 U10687 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n644 ), 
        .Y(n8194) );
  AND2X1 U10688 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[8][6] ), .B(n8901), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n659 )
         );
  INVX1 U10689 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n659 ), 
        .Y(n8195) );
  AND2X1 U10690 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[9][7] ), .B(n8903), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n679 )
         );
  INVX1 U10691 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n679 ), 
        .Y(n8196) );
  AND2X1 U10692 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[10][8] ), .B(n8905), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n698 )
         );
  INVX1 U10693 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n698 ), 
        .Y(n8197) );
  AND2X1 U10694 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[11][9] ), .B(n8907), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n716 )
         );
  INVX1 U10695 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n716 ), 
        .Y(n8198) );
  AND2X1 U10696 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[12][10] ), .B(n8909), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n734 )
         );
  INVX1 U10697 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n734 ), 
        .Y(n8199) );
  AND2X1 U10698 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[13][11] ), .B(n8911), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n752 )
         );
  INVX1 U10699 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n752 ), 
        .Y(n8200) );
  AND2X1 U10700 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][0] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n758 )
         );
  INVX1 U10701 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n758 ), 
        .Y(n8201) );
  AND2X1 U10702 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[14][12] ), .B(n8913), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n770 )
         );
  INVX1 U10703 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n770 ), 
        .Y(n8202) );
  AND2X1 U10704 ( .A(n9466), .B(data_read_reg_1495[14]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n804 )
         );
  INVX1 U10705 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n804 ), 
        .Y(n8203) );
  AND2X1 U10706 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][1] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n810 )
         );
  INVX1 U10707 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n810 ), 
        .Y(n8204) );
  AND2X1 U10708 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[16][13] ), .B(n8915), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n822 )
         );
  INVX1 U10709 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n822 ), 
        .Y(n8205) );
  AND2X1 U10710 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[17][14] ), .B(n8916), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n841 )
         );
  INVX1 U10711 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n841 ), 
        .Y(n8206) );
  AND2X1 U10712 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[18][15] ), .B(n8917), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n859 )
         );
  INVX1 U10713 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n859 ), 
        .Y(n8207) );
  AND2X1 U10714 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 ), 
        .B(data_read_reg_1495[15]), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n892 )
         );
  INVX1 U10715 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n892 ), 
        .Y(n8208) );
  AND2X1 U10716 ( .A(sum_reg_308[31]), .B(n8929), .Y(n2574) );
  INVX1 U10717 ( .A(n2574), .Y(n8209) );
  AND2X1 U10718 ( .A(tmp_7_fu_511_p3[31]), .B(n8965), .Y(n491) );
  INVX1 U10719 ( .A(n491), .Y(n8210) );
  AND2X1 U10720 ( .A(tmp_29_i_fu_752_p2[1]), .B(n8920), .Y(n3173) );
  INVX1 U10721 ( .A(n3173), .Y(n8211) );
  AND2X1 U10722 ( .A(tmp_29_i1_fu_1065_p2[1]), .B(n8922), .Y(n3225) );
  INVX1 U10723 ( .A(n3225), .Y(n8212) );
  AND2X1 U10724 ( .A(sum_reg_308[5]), .B(n8929), .Y(n2678) );
  INVX1 U10725 ( .A(n2678), .Y(n8213) );
  AND2X1 U10726 ( .A(sum_1_reg_376[4]), .B(n8930), .Y(n2424) );
  INVX1 U10727 ( .A(n2424), .Y(n8214) );
  AND2X1 U10728 ( .A(sum_1_reg_376[17]), .B(n8930), .Y(n2476) );
  INVX1 U10729 ( .A(n2476), .Y(n8215) );
  AND2X1 U10730 ( .A(tmp_29_i_fu_752_p2[31]), .B(n8920), .Y(n3160) );
  INVX1 U10731 ( .A(n3160), .Y(n8216) );
  OR2X1 U10732 ( .A(recentVBools_sum[30]), .B(n8830), .Y(n8850) );
  AND2X1 U10733 ( .A(tmp_29_i1_fu_1065_p2[31]), .B(n8922), .Y(n3212) );
  INVX1 U10734 ( .A(n3212), .Y(n8217) );
  OR2X1 U10735 ( .A(recentABools_sum[30]), .B(n8829), .Y(n8851) );
  INVX1 U10736 ( .A(n4054), .Y(n8218) );
  AND2X1 U10737 ( .A(\toReturn_8_reg_1755[0] ), .B(n10535), .Y(n2048) );
  INVX1 U10738 ( .A(n2048), .Y(n8219) );
  BUFX2 U10739 ( .A(n2049), .Y(n8220) );
  INVX1 U10740 ( .A(n3783), .Y(n8221) );
  AND2X1 U10741 ( .A(\toReturn_6_reg_1660[0] ), .B(n10057), .Y(n1513) );
  INVX1 U10742 ( .A(n1513), .Y(n8222) );
  BUFX2 U10743 ( .A(n1514), .Y(n8223) );
  INVX1 U10744 ( .A(n4616), .Y(n8224) );
  AND2X1 U10745 ( .A(ACaptureThresh_loc_reg_288[18]), .B(n8971), .Y(n3026) );
  INVX1 U10746 ( .A(n3026), .Y(n8225) );
  BUFX2 U10747 ( .A(n3025), .Y(n8226) );
  INVX1 U10748 ( .A(n4569), .Y(n8227) );
  AND2X1 U10749 ( .A(VCaptureThresh_loc_reg_298[1]), .B(n8971), .Y(n2932) );
  INVX1 U10750 ( .A(n2932), .Y(n8228) );
  BUFX2 U10751 ( .A(n2931), .Y(n8229) );
  INVX1 U10752 ( .A(n4556), .Y(n8230) );
  AND2X1 U10753 ( .A(VCaptureThresh_loc_reg_298[14]), .B(n8970), .Y(n2906) );
  INVX1 U10754 ( .A(n2906), .Y(n8231) );
  BUFX2 U10755 ( .A(n2905), .Y(n8232) );
  INVX1 U10756 ( .A(n4540), .Y(n8233) );
  AND2X1 U10757 ( .A(VCaptureThresh_loc_reg_298[30]), .B(n8969), .Y(n2874) );
  INVX1 U10758 ( .A(n2874), .Y(n8234) );
  BUFX2 U10759 ( .A(n2873), .Y(n8235) );
  OR2X1 U10760 ( .A(VbeatFallDelay_new_1_reg_342[22]), .B(
        VbeatFallDelay_new_1_reg_342[21]), .Y(n11904) );
  INVX1 U10761 ( .A(n11904), .Y(n8236) );
  AND2X1 U10762 ( .A(tmp_6_reg_1538[13]), .B(n9586), .Y(n11930) );
  INVX1 U10763 ( .A(n11930), .Y(n8237) );
  AND2X1 U10764 ( .A(tmp_7_reg_1544[13]), .B(n9693), .Y(n12019) );
  INVX1 U10765 ( .A(n12019), .Y(n8238) );
  AND2X1 U10766 ( .A(VbeatDelay_new_1_reg_326[13]), .B(n10401), .Y(n11822) );
  INVX1 U10767 ( .A(n11822), .Y(n8239) );
  OR2X1 U10768 ( .A(p_tmp_i_reg_1556[22]), .B(p_tmp_i_reg_1556[21]), .Y(n11244) );
  INVX1 U10769 ( .A(n11244), .Y(n8240) );
  OR2X1 U10770 ( .A(CircularBuffer_head_i_read_ass_reg_1624[7]), .B(n11362), 
        .Y(n11364) );
  INVX1 U10771 ( .A(n11364), .Y(n8241) );
  AND2X1 U10772 ( .A(CircularBuffer_head_i_read_ass_reg_1624[7]), .B(n11362), 
        .Y(n11363) );
  INVX1 U10773 ( .A(n11363), .Y(n8242) );
  OR2X1 U10774 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[7]), .B(n11414), 
        .Y(n11416) );
  INVX1 U10775 ( .A(n11416), .Y(n8243) );
  AND2X1 U10776 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[7]), .B(n11414), 
        .Y(n11415) );
  INVX1 U10777 ( .A(n11415), .Y(n8244) );
  BUFX2 U10778 ( .A(n11952), .Y(n8245) );
  BUFX2 U10779 ( .A(n12041), .Y(n8246) );
  BUFX2 U10780 ( .A(n11120), .Y(n8247) );
  BUFX2 U10781 ( .A(n11835), .Y(n8248) );
  BUFX2 U10782 ( .A(n11832), .Y(n8249) );
  OR2X1 U10783 ( .A(tmp_38_i_reg_1550[20]), .B(tmp_38_i_reg_1550[1]), .Y(n1664) );
  INVX1 U10784 ( .A(n1664), .Y(n8250) );
  OR2X1 U10785 ( .A(CircularBuffer_len_read_assign_1_reg_1616[9]), .B(
        CircularBuffer_len_read_assign_1_reg_1616[8]), .Y(n1504) );
  INVX1 U10786 ( .A(n1504), .Y(n8251) );
  OR2X1 U10787 ( .A(CircularBuffer_len_read_assign_3_reg_1711[9]), .B(
        CircularBuffer_len_read_assign_3_reg_1711[8]), .Y(n869) );
  INVX1 U10788 ( .A(n869), .Y(n8252) );
  OR2X1 U10789 ( .A(p_tmp_i_fu_587_p3[10]), .B(n9886), .Y(n1940) );
  INVX1 U10790 ( .A(n1940), .Y(n8253) );
  OR2X1 U10791 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[9]), .B(
        CircularBuffer_head_i_read_ass_fu_797_p3[8]), .Y(n1819) );
  INVX1 U10792 ( .A(n1819), .Y(n8254) );
  OR2X1 U10793 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[20]), .B(
        CircularBuffer_head_i_read_ass_fu_797_p3[19]), .Y(n1809) );
  INVX1 U10794 ( .A(n1809), .Y(n8255) );
  OR2X1 U10795 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[9]), .B(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[8]), .Y(n1263) );
  INVX1 U10796 ( .A(n1263), .Y(n8256) );
  OR2X1 U10797 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[20]), .B(
        CircularBuffer_head_i_read_ass_1_fu_1110_p3[19]), .Y(n1245) );
  INVX1 U10798 ( .A(n1245), .Y(n8257) );
  OR2X1 U10799 ( .A(tmp_38_i_reg_1550[23]), .B(tmp_38_i_reg_1550[22]), .Y(
        n2059) );
  INVX1 U10800 ( .A(n2059), .Y(n8258) );
  OR2X1 U10801 ( .A(tmp_38_i_reg_1550[9]), .B(tmp_38_i_reg_1550[8]), .Y(n2068)
         );
  INVX1 U10802 ( .A(n2068), .Y(n8259) );
  OR2X1 U10803 ( .A(recentVBools_len[20]), .B(recentVBools_len[19]), .Y(n3193)
         );
  INVX1 U10804 ( .A(n3193), .Y(n8260) );
  OR2X1 U10805 ( .A(recentVBools_len[9]), .B(recentVBools_len[8]), .Y(n3202)
         );
  INVX1 U10806 ( .A(n3202), .Y(n8261) );
  OR2X1 U10807 ( .A(recentABools_len[20]), .B(recentABools_len[19]), .Y(n3245)
         );
  INVX1 U10808 ( .A(n3245), .Y(n8262) );
  OR2X1 U10809 ( .A(recentABools_len[9]), .B(recentABools_len[8]), .Y(n3254)
         );
  INVX1 U10810 ( .A(n3254), .Y(n8263) );
  OR2X1 U10811 ( .A(tmp_38_i_reg_1550[3]), .B(tmp_38_i_reg_1550[31]), .Y(n1685) );
  INVX1 U10812 ( .A(n1685), .Y(n8264) );
  OR2X1 U10813 ( .A(AbeatDelay_new_reg_394[4]), .B(AbeatDelay_new_reg_394[3]), 
        .Y(n298) );
  INVX1 U10814 ( .A(n298), .Y(n8265) );
  OR2X1 U10815 ( .A(n8918), .B(\Decision_AXILiteS_s_axi_U/n315 ), .Y(
        \Decision_AXILiteS_s_axi_U/n629 ) );
  INVX1 U10816 ( .A(\Decision_AXILiteS_s_axi_U/n629 ), .Y(n8266) );
  INVX1 U10817 ( .A(\Decision_AXILiteS_s_axi_U/n332 ), .Y(n8267) );
  BUFX2 U10818 ( .A(\Decision_AXILiteS_s_axi_U/n333 ), .Y(n8268) );
  AND2X1 U10819 ( .A(n9920), .B(n9919), .Y(n1665) );
  INVX1 U10820 ( .A(n1665), .Y(n8269) );
  AND2X1 U10821 ( .A(n10104), .B(n10105), .Y(n1508) );
  INVX1 U10822 ( .A(n1508), .Y(n8270) );
  AND2X1 U10823 ( .A(n10599), .B(n10600), .Y(n873) );
  INVX1 U10824 ( .A(n873), .Y(n8271) );
  AND2X1 U10825 ( .A(ap_CS_fsm[5]), .B(n10139), .Y(n1552) );
  INVX1 U10826 ( .A(n1552), .Y(n8272) );
  AND2X1 U10827 ( .A(ap_CS_fsm[10]), .B(n10634), .Y(n830) );
  INVX1 U10828 ( .A(n830), .Y(n8273) );
  BUFX2 U10829 ( .A(n1476), .Y(n8274) );
  OR2X1 U10830 ( .A(CircularBuffer_len_read_assign_1_reg_1616[23]), .B(
        CircularBuffer_len_read_assign_1_reg_1616[22]), .Y(n1485) );
  INVX1 U10831 ( .A(n1485), .Y(n8275) );
  BUFX2 U10832 ( .A(n841), .Y(n8276) );
  OR2X1 U10833 ( .A(CircularBuffer_len_read_assign_3_reg_1711[23]), .B(
        CircularBuffer_len_read_assign_3_reg_1711[22]), .Y(n850) );
  INVX1 U10834 ( .A(n850), .Y(n8277) );
  AND2X1 U10835 ( .A(vflip[1]), .B(vflip[0]), .Y(n433) );
  INVX1 U10836 ( .A(n433), .Y(n8278) );
  AND2X1 U10837 ( .A(aflip[1]), .B(aflip[0]), .Y(n475) );
  INVX1 U10838 ( .A(n475), .Y(n8279) );
  AND2X1 U10839 ( .A(n10142), .B(n10143), .Y(n1535) );
  INVX1 U10840 ( .A(n1535), .Y(n8280) );
  AND2X1 U10841 ( .A(n10637), .B(n10638), .Y(n813) );
  INVX1 U10842 ( .A(n813), .Y(n8281) );
  AND2X1 U10843 ( .A(n10737), .B(n10681), .Y(n299) );
  INVX1 U10844 ( .A(n299), .Y(n8282) );
  AND2X1 U10845 ( .A(n10136), .B(n10137), .Y(n3203) );
  INVX1 U10846 ( .A(n3203), .Y(n8283) );
  AND2X1 U10847 ( .A(n10631), .B(n10632), .Y(n3255) );
  INVX1 U10848 ( .A(n3255), .Y(n8284) );
  AND2X1 U10849 ( .A(n9830), .B(n9902), .Y(n2069) );
  INVX1 U10850 ( .A(n2069), .Y(n8285) );
  BUFX2 U10851 ( .A(n1540), .Y(n8286) );
  OR2X1 U10852 ( .A(CircularBuffer_len_write_assig_reg_1634[19]), .B(
        CircularBuffer_len_write_assig_reg_1634[18]), .Y(n1543) );
  INVX1 U10853 ( .A(n1543), .Y(n8287) );
  BUFX2 U10854 ( .A(n818), .Y(n8288) );
  OR2X1 U10855 ( .A(CircularBuffer_len_write_assig_2_reg_1729[19]), .B(
        CircularBuffer_len_write_assig_2_reg_1729[18]), .Y(n821) );
  INVX1 U10856 ( .A(n821), .Y(n8289) );
  AND2X1 U10857 ( .A(n9860), .B(n8659), .Y(n1948) );
  INVX1 U10858 ( .A(n1948), .Y(n8290) );
  BUFX2 U10859 ( .A(n1946), .Y(n8291) );
  AND2X1 U10860 ( .A(n8657), .B(n8934), .Y(n2403) );
  INVX1 U10861 ( .A(n2403), .Y(n8292) );
  AND2X1 U10862 ( .A(n8656), .B(n8927), .Y(n2864) );
  INVX1 U10863 ( .A(n2864), .Y(n8293) );
  AND2X1 U10864 ( .A(n367), .B(n8968), .Y(N472) );
  INVX1 U10865 ( .A(N472), .Y(n8294) );
  AND2X1 U10866 ( .A(n11228), .B(n10071), .Y(n11229) );
  INVX1 U10867 ( .A(n11229), .Y(n8295) );
  AND2X1 U10868 ( .A(n11198), .B(n10536), .Y(n11199) );
  INVX1 U10869 ( .A(n11199), .Y(n8296) );
  AND2X1 U10870 ( .A(n11214), .B(n10073), .Y(n11225) );
  INVX1 U10871 ( .A(n11225), .Y(n8297) );
  AND2X1 U10872 ( .A(n11184), .B(n10538), .Y(n11195) );
  INVX1 U10873 ( .A(n11195), .Y(n8298) );
  AND2X1 U10874 ( .A(n9899), .B(n9900), .Y(n11235) );
  INVX1 U10875 ( .A(n11235), .Y(n8299) );
  AND2X1 U10876 ( .A(N512), .B(n8996), .Y(n1646) );
  AND2X1 U10877 ( .A(N497), .B(n9019), .Y(n970) );
  AND2X1 U10878 ( .A(recentdatapoints_len_load_op_fu_556_p2[14]), .B(n8972), 
        .Y(n1836) );
  INVX1 U10879 ( .A(n1836), .Y(n8300) );
  AND2X1 U10880 ( .A(recentdatapoints_len_load_op_fu_556_p2[27]), .B(n8972), 
        .Y(n1854) );
  INVX1 U10881 ( .A(n1854), .Y(n8301) );
  AND2X1 U10882 ( .A(recentdatapoints_len_load_op_fu_556_p2[31]), .B(n8972), 
        .Y(n1859) );
  INVX1 U10883 ( .A(n1859), .Y(n8302) );
  AND2X1 U10884 ( .A(n5965), .B(ap_CS_fsm[12]), .Y(n2155) );
  INVX1 U10885 ( .A(n2155), .Y(n8303) );
  AND2X1 U10886 ( .A(ap_CS_fsm[0]), .B(n10889), .Y(n2154) );
  INVX1 U10887 ( .A(n2154), .Y(n8304) );
  AND2X1 U10888 ( .A(n9935), .B(tmp_33_i_fu_786_p2[1]), .Y(n1695) );
  INVX1 U10889 ( .A(n1695), .Y(n8305) );
  AND2X1 U10890 ( .A(n10243), .B(tmp_33_i1_fu_1099_p2[1]), .Y(n1212) );
  INVX1 U10891 ( .A(n1212), .Y(n8306) );
  BUFX2 U10892 ( .A(n11105), .Y(n8307) );
  OR2X1 U10893 ( .A(AbeatDelay_new_reg_394[10]), .B(AbeatDelay_new_reg_394[11]), .Y(n11062) );
  INVX1 U10894 ( .A(n11062), .Y(n8308) );
  AND2X1 U10895 ( .A(v_thresh[15]), .B(n9535), .Y(n12223) );
  INVX1 U10896 ( .A(n12223), .Y(n8309) );
  AND2X1 U10897 ( .A(v_thresh[11]), .B(n9534), .Y(n12217) );
  INVX1 U10898 ( .A(n12217), .Y(n8310) );
  AND2X1 U10899 ( .A(v_thresh[3]), .B(n9537), .Y(n12202) );
  INVX1 U10900 ( .A(n12202), .Y(n8311) );
  AND2X1 U10901 ( .A(v_thresh[7]), .B(n9538), .Y(n12207) );
  INVX1 U10902 ( .A(n12207), .Y(n8312) );
  AND2X1 U10903 ( .A(a_thresh[11]), .B(n9475), .Y(n11584) );
  INVX1 U10904 ( .A(n11584), .Y(n8313) );
  AND2X1 U10905 ( .A(a_thresh[3]), .B(n9482), .Y(n11569) );
  INVX1 U10906 ( .A(n11569), .Y(n8314) );
  AND2X1 U10907 ( .A(a_thresh[7]), .B(n9485), .Y(n11574) );
  INVX1 U10908 ( .A(n11574), .Y(n8315) );
  AND2X1 U10909 ( .A(ACaptureThresh_loc_reg_288[27]), .B(n10770), .Y(n11967)
         );
  INVX1 U10910 ( .A(n11967), .Y(n8316) );
  AND2X1 U10911 ( .A(ACaptureThresh_loc_reg_288[15]), .B(n10758), .Y(n11927)
         );
  INVX1 U10912 ( .A(n11927), .Y(n8317) );
  AND2X1 U10913 ( .A(ACaptureThresh_loc_reg_288[11]), .B(n10754), .Y(n11921)
         );
  INVX1 U10914 ( .A(n11921), .Y(n8318) );
  AND2X1 U10915 ( .A(VCaptureThresh_loc_reg_298[27]), .B(n10804), .Y(n12056)
         );
  INVX1 U10916 ( .A(n12056), .Y(n8319) );
  AND2X1 U10917 ( .A(VCaptureThresh_loc_reg_298[15]), .B(n10792), .Y(n12016)
         );
  INVX1 U10918 ( .A(n12016), .Y(n8320) );
  AND2X1 U10919 ( .A(VCaptureThresh_loc_reg_298[11]), .B(n10788), .Y(n12010)
         );
  INVX1 U10920 ( .A(n12010), .Y(n8321) );
  AND2X1 U10921 ( .A(VCaptureThresh_loc_reg_298[28]), .B(n10069), .Y(n11512)
         );
  INVX1 U10922 ( .A(n11512), .Y(n8322) );
  AND2X1 U10923 ( .A(n2862), .B(n9765), .Y(n12152) );
  INVX1 U10924 ( .A(n12152), .Y(n8323) );
  AND2X1 U10925 ( .A(n2401), .B(n9646), .Y(n11688) );
  INVX1 U10926 ( .A(n11688), .Y(n8324) );
  AND2X1 U10927 ( .A(VbeatDelay_new_1_reg_326[31]), .B(n10741), .Y(n11142) );
  INVX1 U10928 ( .A(n11142), .Y(n8325) );
  AND2X1 U10929 ( .A(VCaptureThresh_loc_reg_298[16]), .B(n10066), .Y(n11472)
         );
  INVX1 U10930 ( .A(n11472), .Y(n8326) );
  AND2X1 U10931 ( .A(VCaptureThresh_loc_reg_298[12]), .B(n10065), .Y(n11466)
         );
  INVX1 U10932 ( .A(n11466), .Y(n8327) );
  AND2X1 U10933 ( .A(VbeatFallDelay_new_1_reg_342[27]), .B(n10523), .Y(n11859)
         );
  INVX1 U10934 ( .A(n11859), .Y(n8328) );
  AND2X1 U10935 ( .A(VbeatFallDelay_new_1_reg_342[15]), .B(n10491), .Y(n11819)
         );
  INVX1 U10936 ( .A(n11819), .Y(n8329) );
  AND2X1 U10937 ( .A(VbeatFallDelay_new_1_reg_342[11]), .B(n10480), .Y(n11813)
         );
  INVX1 U10938 ( .A(n11813), .Y(n8330) );
  AND2X1 U10939 ( .A(ACaptureThresh_loc_reg_288[28]), .B(n9332), .Y(n11770) );
  INVX1 U10940 ( .A(n11770), .Y(n8331) );
  AND2X1 U10941 ( .A(ACaptureThresh_loc_reg_288[16]), .B(n9356), .Y(n11730) );
  INVX1 U10942 ( .A(n11730), .Y(n8332) );
  AND2X1 U10943 ( .A(ACaptureThresh_loc_reg_288[12]), .B(n9363), .Y(n11724) );
  INVX1 U10944 ( .A(n11724), .Y(n8333) );
  AND2X1 U10945 ( .A(ACaptureThresh_loc_reg_288[23]), .B(n10766), .Y(n11991)
         );
  INVX1 U10946 ( .A(n11991), .Y(n8334) );
  AND2X1 U10947 ( .A(ACaptureThresh_loc_reg_288[19]), .B(n10762), .Y(n11984)
         );
  INVX1 U10948 ( .A(n11984), .Y(n8335) );
  AND2X1 U10949 ( .A(VCaptureThresh_loc_reg_298[23]), .B(n10800), .Y(n12080)
         );
  INVX1 U10950 ( .A(n12080), .Y(n8336) );
  AND2X1 U10951 ( .A(VCaptureThresh_loc_reg_298[19]), .B(n10796), .Y(n12073)
         );
  INVX1 U10952 ( .A(n12073), .Y(n8337) );
  AND2X1 U10953 ( .A(VCaptureThresh_loc_reg_298[20]), .B(n10067), .Y(n11529)
         );
  INVX1 U10954 ( .A(n11529), .Y(n8338) );
  AND2X1 U10955 ( .A(VCaptureThresh_loc_reg_298[8]), .B(n10063), .Y(n11492) );
  INVX1 U10956 ( .A(n11492), .Y(n8339) );
  AND2X1 U10957 ( .A(VbeatFallDelay_new_1_reg_342[23]), .B(n10512), .Y(n11883)
         );
  INVX1 U10958 ( .A(n11883), .Y(n8340) );
  AND2X1 U10959 ( .A(VbeatFallDelay_new_1_reg_342[19]), .B(n10501), .Y(n11876)
         );
  INVX1 U10960 ( .A(n11876), .Y(n8341) );
  AND2X1 U10961 ( .A(ACaptureThresh_loc_reg_288[24]), .B(n9340), .Y(n11794) );
  INVX1 U10962 ( .A(n11794), .Y(n8342) );
  AND2X1 U10963 ( .A(ACaptureThresh_loc_reg_288[20]), .B(n9347), .Y(n11787) );
  INVX1 U10964 ( .A(n11787), .Y(n8343) );
  AND2X1 U10965 ( .A(ACaptureThresh_loc_reg_288[7]), .B(n10750), .Y(n11947) );
  INVX1 U10966 ( .A(n11947), .Y(n8344) );
  AND2X1 U10967 ( .A(VCaptureThresh_loc_reg_298[7]), .B(n10784), .Y(n12036) );
  INVX1 U10968 ( .A(n12036), .Y(n8345) );
  AND2X1 U10969 ( .A(VCaptureThresh_loc_reg_298[24]), .B(n10068), .Y(n11536)
         );
  INVX1 U10970 ( .A(n11536), .Y(n8346) );
  AND2X1 U10971 ( .A(VbeatFallDelay_new_1_reg_342[3]), .B(n10459), .Y(n11836)
         );
  INVX1 U10972 ( .A(n11836), .Y(n8347) );
  AND2X1 U10973 ( .A(VbeatFallDelay_new_1_reg_342[7]), .B(n10468), .Y(n11839)
         );
  INVX1 U10974 ( .A(n11839), .Y(n8348) );
  AND2X1 U10975 ( .A(ACaptureThresh_loc_reg_288[4]), .B(n9377), .Y(n11747) );
  INVX1 U10976 ( .A(n11747), .Y(n8349) );
  AND2X1 U10977 ( .A(ACaptureThresh_loc_reg_288[8]), .B(n9371), .Y(n11750) );
  INVX1 U10978 ( .A(n11750), .Y(n8350) );
  AND2X1 U10979 ( .A(VCaptureThresh_loc_reg_298[3]), .B(n10072), .Y(n12122) );
  INVX1 U10980 ( .A(n12122), .Y(n8351) );
  AND2X1 U10981 ( .A(ACaptureThresh_loc_reg_288[3]), .B(n10537), .Y(n11658) );
  INVX1 U10982 ( .A(n11658), .Y(n8352) );
  AND2X1 U10983 ( .A(VCaptureThresh_loc_reg_298[4]), .B(n10062), .Y(n11489) );
  INVX1 U10984 ( .A(n11489), .Y(n8353) );
  AND2X1 U10985 ( .A(\Decision_AXILiteS_s_axi_U/wstate[1] ), .B(n10901), .Y(
        s_axi_AXILiteS_BVALID) );
  INVX1 U10986 ( .A(s_axi_AXILiteS_BVALID), .Y(n8354) );
  AND2X1 U10987 ( .A(n8978), .B(n9013), .Y(n364) );
  INVX1 U10988 ( .A(n364), .Y(n8355) );
  OR2X1 U10989 ( .A(n9507), .B(p_cast_fu_688_p1[9]), .Y(n12236) );
  INVX1 U10990 ( .A(n12236), .Y(n8356) );
  OR2X1 U10991 ( .A(n9771), .B(p_1_cast_fu_1031_p1[9]), .Y(n11603) );
  INVX1 U10992 ( .A(n11603), .Y(n8357) );
  OR2X1 U10993 ( .A(n9573), .B(tmp_6_reg_1538[9]), .Y(n11938) );
  INVX1 U10994 ( .A(n11938), .Y(n8358) );
  OR2X1 U10995 ( .A(n9677), .B(tmp_7_reg_1544[9]), .Y(n12027) );
  INVX1 U10996 ( .A(n12027), .Y(n8359) );
  OR2X1 U10997 ( .A(n10390), .B(VbeatDelay_new_1_reg_326[9]), .Y(n11830) );
  INVX1 U10998 ( .A(n11830), .Y(n8360) );
  OR2X1 U10999 ( .A(n9579), .B(sum_1_phi_fu_379_p4[9]), .Y(n11741) );
  INVX1 U11000 ( .A(n11741), .Y(n8361) );
  OR2X1 U11001 ( .A(n9683), .B(sum_phi_fu_311_p4[9]), .Y(n11483) );
  INVX1 U11002 ( .A(n11483), .Y(n8362) );
  BUFX2 U11003 ( .A(n11358), .Y(n8363) );
  BUFX2 U11004 ( .A(n11356), .Y(n8364) );
  BUFX2 U11005 ( .A(n11355), .Y(n8365) );
  BUFX2 U11006 ( .A(n11462), .Y(n8366) );
  BUFX2 U11007 ( .A(n11460), .Y(n8367) );
  BUFX2 U11008 ( .A(n11459), .Y(n8368) );
  BUFX2 U11009 ( .A(n11309), .Y(n8369) );
  BUFX2 U11010 ( .A(n11257), .Y(n8370) );
  BUFX2 U11011 ( .A(n12253), .Y(n8371) );
  BUFX2 U11012 ( .A(n11620), .Y(n8372) );
  BUFX2 U11013 ( .A(n11983), .Y(n8373) );
  BUFX2 U11014 ( .A(n12072), .Y(n8374) );
  BUFX2 U11015 ( .A(n11875), .Y(n8375) );
  BUFX2 U11016 ( .A(n11528), .Y(n8376) );
  BUFX2 U11017 ( .A(n11786), .Y(n8377) );
  AND2X1 U11018 ( .A(N495), .B(ap_CS_fsm[7]), .Y(n2567) );
  INVX1 U11019 ( .A(n2567), .Y(n8378) );
  INVX1 U11020 ( .A(n2018), .Y(n8379) );
  BUFX2 U11021 ( .A(n2028), .Y(n8380) );
  BUFX2 U11022 ( .A(n2029), .Y(n8381) );
  INVX1 U11023 ( .A(\Decision_AXILiteS_s_axi_U/n576 ), .Y(n8382) );
  BUFX2 U11024 ( .A(\Decision_AXILiteS_s_axi_U/n319 ), .Y(n8383) );
  AND2X1 U11025 ( .A(n11246), .B(n9897), .Y(n11254) );
  INVX1 U11026 ( .A(n11254), .Y(n8384) );
  INVX1 U11027 ( .A(n11226), .Y(n8385) );
  INVX1 U11028 ( .A(n11196), .Y(n8386) );
  AND2X1 U11029 ( .A(recentdatapoints_data_q0[12]), .B(n8868), .Y(n423) );
  INVX1 U11030 ( .A(n423), .Y(n8387) );
  AND2X1 U11031 ( .A(n9281), .B(ap_rst_n), .Y(\Decision_AXILiteS_s_axi_U/n599 ) );
  INVX1 U11032 ( .A(\Decision_AXILiteS_s_axi_U/n599 ), .Y(n8388) );
  AND2X1 U11033 ( .A(s_axi_AXILiteS_WDATA[0]), .B(
        \Decision_AXILiteS_s_axi_U/n617 ), .Y(\Decision_AXILiteS_s_axi_U/n564 ) );
  INVX1 U11034 ( .A(\Decision_AXILiteS_s_axi_U/n564 ), .Y(n8389) );
  AND2X1 U11035 ( .A(recentdatapoints_data_q0[0]), .B(n8869), .Y(n429) );
  INVX1 U11036 ( .A(n429), .Y(n8390) );
  AND2X1 U11037 ( .A(n10075), .B(n3151), .Y(n2794) );
  INVX1 U11038 ( .A(n2794), .Y(n8391) );
  AND2X1 U11039 ( .A(n10540), .B(n3149), .Y(n2301) );
  INVX1 U11040 ( .A(n2301), .Y(n8392) );
  INVX1 U11041 ( .A(\toReturn_1_fu_1395_p3[7] ), .Y(n8393) );
  BUFX2 U11042 ( .A(n305), .Y(n8394) );
  BUFX2 U11043 ( .A(n306), .Y(n8395) );
  BUFX2 U11044 ( .A(n2199), .Y(n8396) );
  OR2X1 U11045 ( .A(n9013), .B(n8975), .Y(n350) );
  INVX1 U11046 ( .A(n350), .Y(n8397) );
  AND2X1 U11047 ( .A(CircularBuffer_len_read_assign_fu_772_p2[11]), .B(n3151), 
        .Y(n2772) );
  INVX1 U11048 ( .A(n2772), .Y(n8398) );
  AND2X1 U11049 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[11]), .B(
        n3149), .Y(n2279) );
  INVX1 U11050 ( .A(n2279), .Y(n8399) );
  AND2X1 U11051 ( .A(CircularBuffer_len_read_assign_fu_772_p2[23]), .B(n8919), 
        .Y(n2748) );
  INVX1 U11052 ( .A(n2748), .Y(n8400) );
  AND2X1 U11053 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[23]), .B(
        n8921), .Y(n2255) );
  INVX1 U11054 ( .A(n2255), .Y(n8401) );
  INVX1 U11055 ( .A(recentABools_data_address0[3]), .Y(n8402) );
  BUFX2 U11056 ( .A(n388), .Y(n8403) );
  BUFX2 U11057 ( .A(n389), .Y(n8404) );
  BUFX2 U11058 ( .A(n2193), .Y(n8405) );
  AND2X1 U11059 ( .A(CircularBuffer_len_read_assign_fu_772_p2[8]), .B(n8919), 
        .Y(n2778) );
  INVX1 U11060 ( .A(n2778), .Y(n8406) );
  AND2X1 U11061 ( .A(CircularBuffer_len_read_assign_2_fu_1085_p2[8]), .B(n3149), .Y(n2285) );
  INVX1 U11062 ( .A(n2285), .Y(n8407) );
  AND2X1 U11063 ( .A(\tmp_i3_reg_1674[0] ), .B(recentdatapoints_data_q0[15]), 
        .Y(n440) );
  INVX1 U11064 ( .A(n440), .Y(n8408) );
  AND2X1 U11065 ( .A(\Decision_AXILiteS_s_axi_U/n351 ), .B(
        \Decision_AXILiteS_s_axi_U/n352 ), .Y(\Decision_AXILiteS_s_axi_U/n343 ) );
  INVX1 U11066 ( .A(\Decision_AXILiteS_s_axi_U/n343 ), .Y(n8409) );
  AND2X1 U11067 ( .A(n8881), .B(\Decision_AXILiteS_s_axi_U/n384 ), .Y(
        \Decision_AXILiteS_s_axi_U/n375 ) );
  INVX1 U11068 ( .A(\Decision_AXILiteS_s_axi_U/n375 ), .Y(n8410) );
  INVX1 U11069 ( .A(\Decision_AXILiteS_s_axi_U/n462 ), .Y(n8411) );
  BUFX2 U11070 ( .A(\Decision_AXILiteS_s_axi_U/n470 ), .Y(n8412) );
  INVX1 U11071 ( .A(recentVBools_data_address0[2]), .Y(n8413) );
  BUFX2 U11072 ( .A(n376), .Y(n8414) );
  BUFX2 U11073 ( .A(n377), .Y(n8415) );
  BUFX2 U11074 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n42 ), .Y(n8416) );
  AND2X1 U11075 ( .A(\Decision_AXILiteS_s_axi_U/n353 ), .B(
        \Decision_AXILiteS_s_axi_U/n429 ), .Y(\Decision_AXILiteS_s_axi_U/n440 ) );
  INVX1 U11076 ( .A(\Decision_AXILiteS_s_axi_U/n440 ), .Y(n8417) );
  AND2X1 U11077 ( .A(\Decision_AXILiteS_s_axi_U/n397 ), .B(n8882), .Y(
        \Decision_AXILiteS_s_axi_U/n493 ) );
  INVX1 U11078 ( .A(\Decision_AXILiteS_s_axi_U/n493 ), .Y(n8418) );
  AND2X1 U11079 ( .A(\Decision_AXILiteS_s_axi_U/n385 ), .B(
        \Decision_AXILiteS_s_axi_U/n533 ), .Y(\Decision_AXILiteS_s_axi_U/n523 ) );
  INVX1 U11080 ( .A(\Decision_AXILiteS_s_axi_U/n523 ), .Y(n8419) );
  INVX1 U11081 ( .A(n8292), .Y(n8890) );
  INVX1 U11082 ( .A(n8293), .Y(n8893) );
  INVX1 U11083 ( .A(n8933), .Y(n8932) );
  INVX1 U11084 ( .A(n8926), .Y(n8925) );
  INVX1 U11085 ( .A(n8892), .Y(n8891) );
  INVX1 U11086 ( .A(n8895), .Y(n8894) );
  INVX1 U11087 ( .A(n2701), .Y(n8926) );
  INVX1 U11088 ( .A(n2241), .Y(n8933) );
  INVX1 U11089 ( .A(n970), .Y(n8892) );
  INVX1 U11090 ( .A(n1646), .Y(n8895) );
  INVX1 U11091 ( .A(n8928), .Y(n8927) );
  INVX1 U11092 ( .A(n8935), .Y(n8934) );
  BUFX2 U11093 ( .A(n9273), .Y(n9070) );
  BUFX2 U11094 ( .A(n9273), .Y(n9071) );
  BUFX2 U11095 ( .A(n9273), .Y(n9072) );
  BUFX2 U11096 ( .A(n9272), .Y(n9073) );
  BUFX2 U11097 ( .A(n9272), .Y(n9074) );
  BUFX2 U11098 ( .A(n9272), .Y(n9075) );
  BUFX2 U11099 ( .A(n9271), .Y(n9076) );
  BUFX2 U11100 ( .A(n9271), .Y(n9077) );
  BUFX2 U11101 ( .A(n9271), .Y(n9078) );
  BUFX2 U11102 ( .A(n9270), .Y(n9079) );
  BUFX2 U11103 ( .A(n9270), .Y(n9080) );
  BUFX2 U11104 ( .A(n9270), .Y(n9081) );
  BUFX2 U11105 ( .A(n9269), .Y(n9082) );
  BUFX2 U11106 ( .A(n9269), .Y(n9083) );
  BUFX2 U11107 ( .A(n9269), .Y(n9084) );
  BUFX2 U11108 ( .A(n9268), .Y(n9085) );
  BUFX2 U11109 ( .A(n9268), .Y(n9086) );
  BUFX2 U11110 ( .A(n9268), .Y(n9087) );
  BUFX2 U11111 ( .A(n9267), .Y(n9088) );
  BUFX2 U11112 ( .A(n9267), .Y(n9089) );
  BUFX2 U11113 ( .A(n9267), .Y(n9090) );
  BUFX2 U11114 ( .A(n9266), .Y(n9091) );
  BUFX2 U11115 ( .A(n9266), .Y(n9092) );
  BUFX2 U11116 ( .A(n9266), .Y(n9093) );
  BUFX2 U11117 ( .A(n9265), .Y(n9094) );
  BUFX2 U11118 ( .A(n9265), .Y(n9095) );
  BUFX2 U11119 ( .A(n9265), .Y(n9096) );
  BUFX2 U11120 ( .A(n9264), .Y(n9097) );
  BUFX2 U11121 ( .A(n9264), .Y(n9098) );
  BUFX2 U11122 ( .A(n9264), .Y(n9099) );
  BUFX2 U11123 ( .A(n9263), .Y(n9100) );
  BUFX2 U11124 ( .A(n9263), .Y(n9101) );
  BUFX2 U11125 ( .A(n9263), .Y(n9102) );
  BUFX2 U11126 ( .A(n9262), .Y(n9103) );
  BUFX2 U11127 ( .A(n9262), .Y(n9104) );
  BUFX2 U11128 ( .A(n9262), .Y(n9105) );
  BUFX2 U11129 ( .A(n9261), .Y(n9106) );
  BUFX2 U11130 ( .A(n9261), .Y(n9107) );
  BUFX2 U11131 ( .A(n9261), .Y(n9108) );
  BUFX2 U11132 ( .A(n9260), .Y(n9109) );
  BUFX2 U11133 ( .A(n9260), .Y(n9110) );
  BUFX2 U11134 ( .A(n9260), .Y(n9111) );
  BUFX2 U11135 ( .A(n9259), .Y(n9112) );
  BUFX2 U11136 ( .A(n9259), .Y(n9113) );
  BUFX2 U11137 ( .A(n9259), .Y(n9114) );
  BUFX2 U11138 ( .A(n9258), .Y(n9115) );
  BUFX2 U11139 ( .A(n9258), .Y(n9116) );
  BUFX2 U11140 ( .A(n9258), .Y(n9117) );
  BUFX2 U11141 ( .A(n9257), .Y(n9118) );
  BUFX2 U11142 ( .A(n9257), .Y(n9119) );
  BUFX2 U11143 ( .A(n9257), .Y(n9120) );
  BUFX2 U11144 ( .A(n9256), .Y(n9121) );
  BUFX2 U11145 ( .A(n9256), .Y(n9122) );
  BUFX2 U11146 ( .A(n9256), .Y(n9123) );
  BUFX2 U11147 ( .A(n9255), .Y(n9124) );
  BUFX2 U11148 ( .A(n9255), .Y(n9125) );
  BUFX2 U11149 ( .A(n9255), .Y(n9126) );
  BUFX2 U11150 ( .A(n9254), .Y(n9127) );
  BUFX2 U11151 ( .A(n9254), .Y(n9128) );
  BUFX2 U11152 ( .A(n9254), .Y(n9129) );
  BUFX2 U11153 ( .A(n9253), .Y(n9130) );
  BUFX2 U11154 ( .A(n9253), .Y(n9131) );
  BUFX2 U11155 ( .A(n9253), .Y(n9132) );
  BUFX2 U11156 ( .A(n9252), .Y(n9133) );
  BUFX2 U11157 ( .A(n9252), .Y(n9134) );
  BUFX2 U11158 ( .A(n9252), .Y(n9135) );
  BUFX2 U11159 ( .A(n9251), .Y(n9136) );
  BUFX2 U11160 ( .A(n9251), .Y(n9137) );
  BUFX2 U11161 ( .A(n9251), .Y(n9138) );
  BUFX2 U11162 ( .A(n9250), .Y(n9139) );
  BUFX2 U11163 ( .A(n9250), .Y(n9140) );
  BUFX2 U11164 ( .A(n9250), .Y(n9141) );
  BUFX2 U11165 ( .A(n9249), .Y(n9142) );
  BUFX2 U11166 ( .A(n9249), .Y(n9143) );
  BUFX2 U11167 ( .A(n9249), .Y(n9144) );
  BUFX2 U11168 ( .A(n9248), .Y(n9145) );
  BUFX2 U11169 ( .A(n9248), .Y(n9146) );
  BUFX2 U11170 ( .A(n9248), .Y(n9147) );
  BUFX2 U11171 ( .A(n9247), .Y(n9148) );
  BUFX2 U11172 ( .A(n9247), .Y(n9149) );
  BUFX2 U11173 ( .A(n9247), .Y(n9150) );
  BUFX2 U11174 ( .A(n9246), .Y(n9151) );
  BUFX2 U11175 ( .A(n9246), .Y(n9152) );
  BUFX2 U11176 ( .A(n9246), .Y(n9153) );
  BUFX2 U11177 ( .A(n9245), .Y(n9154) );
  BUFX2 U11178 ( .A(n9245), .Y(n9155) );
  BUFX2 U11179 ( .A(n9245), .Y(n9156) );
  BUFX2 U11180 ( .A(n9244), .Y(n9157) );
  BUFX2 U11181 ( .A(n9244), .Y(n9158) );
  BUFX2 U11182 ( .A(n9244), .Y(n9159) );
  BUFX2 U11183 ( .A(n9243), .Y(n9160) );
  BUFX2 U11184 ( .A(n9243), .Y(n9161) );
  BUFX2 U11185 ( .A(n9243), .Y(n9162) );
  BUFX2 U11186 ( .A(n9242), .Y(n9163) );
  BUFX2 U11187 ( .A(n9242), .Y(n9164) );
  BUFX2 U11188 ( .A(n9242), .Y(n9165) );
  BUFX2 U11189 ( .A(n9241), .Y(n9166) );
  BUFX2 U11190 ( .A(n9241), .Y(n9167) );
  BUFX2 U11191 ( .A(n9241), .Y(n9168) );
  BUFX2 U11192 ( .A(n9240), .Y(n9169) );
  BUFX2 U11193 ( .A(n9240), .Y(n9170) );
  BUFX2 U11194 ( .A(n9240), .Y(n9171) );
  BUFX2 U11195 ( .A(n9239), .Y(n9172) );
  BUFX2 U11196 ( .A(n9239), .Y(n9173) );
  BUFX2 U11197 ( .A(n9239), .Y(n9174) );
  BUFX2 U11198 ( .A(n9238), .Y(n9175) );
  BUFX2 U11199 ( .A(n9238), .Y(n9176) );
  BUFX2 U11200 ( .A(n9238), .Y(n9177) );
  BUFX2 U11201 ( .A(n9237), .Y(n9178) );
  BUFX2 U11202 ( .A(n9237), .Y(n9179) );
  BUFX2 U11203 ( .A(n9237), .Y(n9180) );
  BUFX2 U11204 ( .A(n9236), .Y(n9181) );
  BUFX2 U11205 ( .A(n9236), .Y(n9182) );
  BUFX2 U11206 ( .A(n9236), .Y(n9183) );
  BUFX2 U11207 ( .A(n9235), .Y(n9184) );
  BUFX2 U11208 ( .A(n9235), .Y(n9185) );
  BUFX2 U11209 ( .A(n9235), .Y(n9186) );
  BUFX2 U11210 ( .A(n9234), .Y(n9187) );
  BUFX2 U11211 ( .A(n9234), .Y(n9188) );
  BUFX2 U11212 ( .A(n9234), .Y(n9189) );
  BUFX2 U11213 ( .A(n9233), .Y(n9190) );
  BUFX2 U11214 ( .A(n9233), .Y(n9191) );
  BUFX2 U11215 ( .A(n9233), .Y(n9192) );
  BUFX2 U11216 ( .A(n9232), .Y(n9193) );
  BUFX2 U11217 ( .A(n9232), .Y(n9194) );
  BUFX2 U11218 ( .A(n9232), .Y(n9195) );
  BUFX2 U11219 ( .A(n9231), .Y(n9196) );
  BUFX2 U11220 ( .A(n9231), .Y(n9197) );
  BUFX2 U11221 ( .A(n9231), .Y(n9198) );
  BUFX2 U11222 ( .A(n9230), .Y(n9199) );
  BUFX2 U11223 ( .A(n9230), .Y(n9200) );
  BUFX2 U11224 ( .A(n9230), .Y(n9201) );
  BUFX2 U11225 ( .A(n9229), .Y(n9202) );
  BUFX2 U11226 ( .A(n9229), .Y(n9203) );
  BUFX2 U11227 ( .A(n9229), .Y(n9204) );
  BUFX2 U11228 ( .A(n9228), .Y(n9205) );
  BUFX2 U11229 ( .A(n9228), .Y(n9206) );
  BUFX2 U11230 ( .A(n9228), .Y(n9207) );
  BUFX2 U11231 ( .A(n9227), .Y(n9208) );
  BUFX2 U11232 ( .A(n9227), .Y(n9209) );
  BUFX2 U11233 ( .A(n9227), .Y(n9210) );
  BUFX2 U11234 ( .A(n9226), .Y(n9211) );
  BUFX2 U11235 ( .A(n9226), .Y(n9212) );
  BUFX2 U11236 ( .A(n9226), .Y(n9213) );
  BUFX2 U11237 ( .A(n9225), .Y(n9214) );
  BUFX2 U11238 ( .A(n9225), .Y(n9215) );
  BUFX2 U11239 ( .A(n9225), .Y(n9216) );
  BUFX2 U11240 ( .A(n9224), .Y(n9217) );
  BUFX2 U11241 ( .A(n9224), .Y(n9218) );
  BUFX2 U11242 ( .A(n9224), .Y(n9219) );
  BUFX2 U11243 ( .A(n9223), .Y(n9220) );
  BUFX2 U11244 ( .A(n9223), .Y(n9221) );
  BUFX2 U11245 ( .A(n9223), .Y(n9222) );
  INVX1 U11246 ( .A(n2239), .Y(n8935) );
  INVX1 U11247 ( .A(n2699), .Y(n8928) );
  INVX1 U11248 ( .A(n8420), .Y(n8915) );
  INVX1 U11249 ( .A(n8421), .Y(n8931) );
  INVX1 U11250 ( .A(n8422), .Y(n8924) );
  INVX1 U11251 ( .A(n8960), .Y(n8940) );
  INVX1 U11252 ( .A(n8956), .Y(n8952) );
  INVX1 U11253 ( .A(n8969), .Y(n8963) );
  INVX1 U11254 ( .A(n8970), .Y(n8964) );
  INVX1 U11255 ( .A(n8958), .Y(n8951) );
  INVX1 U11256 ( .A(n8957), .Y(n8941) );
  INVX1 U11257 ( .A(n8960), .Y(n8943) );
  INVX1 U11258 ( .A(n8958), .Y(n8942) );
  INVX1 U11259 ( .A(n8960), .Y(n8944) );
  INVX1 U11260 ( .A(n8956), .Y(n8945) );
  INVX1 U11261 ( .A(n8960), .Y(n8950) );
  INVX1 U11262 ( .A(n8956), .Y(n8949) );
  INVX1 U11263 ( .A(n8959), .Y(n8948) );
  INVX1 U11264 ( .A(n8960), .Y(n8946) );
  INVX1 U11265 ( .A(n8957), .Y(n8947) );
  INVX1 U11266 ( .A(n8969), .Y(n8961) );
  INVX1 U11267 ( .A(n8968), .Y(n8962) );
  INVX1 U11268 ( .A(n8958), .Y(n8939) );
  INVX1 U11269 ( .A(n8958), .Y(n8936) );
  INVX1 U11270 ( .A(n8960), .Y(n8937) );
  INVX1 U11271 ( .A(n8959), .Y(n8938) );
  INVX1 U11272 ( .A(n9014), .Y(n9036) );
  INVX1 U11273 ( .A(n9014), .Y(n9035) );
  INVX1 U11274 ( .A(ap_CS_fsm[9]), .Y(n9032) );
  INVX1 U11275 ( .A(n9014), .Y(n9033) );
  INVX1 U11276 ( .A(ap_CS_fsm[9]), .Y(n9034) );
  INVX1 U11277 ( .A(n9014), .Y(n9031) );
  INVX1 U11278 ( .A(ap_CS_fsm[9]), .Y(n9026) );
  INVX1 U11279 ( .A(n9014), .Y(n9025) );
  INVX1 U11280 ( .A(n9017), .Y(n9024) );
  INVX1 U11281 ( .A(n9014), .Y(n9022) );
  INVX1 U11282 ( .A(ap_CS_fsm[9]), .Y(n9023) );
  INVX1 U11283 ( .A(n9014), .Y(n9027) );
  INVX1 U11284 ( .A(n9014), .Y(n9028) );
  INVX1 U11285 ( .A(ap_CS_fsm[9]), .Y(n9029) );
  INVX1 U11286 ( .A(n9014), .Y(n9030) );
  INVX1 U11287 ( .A(n9014), .Y(n9021) );
  INVX1 U11288 ( .A(n9017), .Y(n9040) );
  BUFX2 U11289 ( .A(n9274), .Y(n9067) );
  BUFX2 U11290 ( .A(n9274), .Y(n9068) );
  BUFX2 U11291 ( .A(n9274), .Y(n9069) );
  AND2X1 U11292 ( .A(ap_rst_n), .B(n8883), .Y(\Decision_AXILiteS_s_axi_U/n579 ) );
  OR2X1 U11293 ( .A(n9005), .B(N512), .Y(n2699) );
  OR2X1 U11294 ( .A(n9031), .B(N497), .Y(n2239) );
  AND2X1 U11295 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n825 ), 
        .B(n8877), .Y(n8420) );
  BUFX2 U11296 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n32 ), 
        .Y(n8864) );
  BUFX2 U11297 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n32 ), 
        .Y(n8865) );
  BUFX2 U11298 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n25 ), 
        .Y(n8860) );
  BUFX2 U11299 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n25 ), 
        .Y(n8861) );
  OR2X1 U11300 ( .A(n9041), .B(n8657), .Y(n8421) );
  OR2X1 U11301 ( .A(n9013), .B(n8656), .Y(n8422) );
  BUFX2 U11302 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n31 ), 
        .Y(n8866) );
  BUFX2 U11303 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n31 ), 
        .Y(n8867) );
  BUFX2 U11304 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n24 ), 
        .Y(n8862) );
  BUFX2 U11305 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n24 ), 
        .Y(n8863) );
  INVX1 U11306 ( .A(n8904), .Y(n8903) );
  INVX1 U11307 ( .A(n8902), .Y(n8901) );
  INVX1 U11308 ( .A(n8912), .Y(n8911) );
  INVX1 U11309 ( .A(n8910), .Y(n8909) );
  INVX1 U11310 ( .A(n8914), .Y(n8913) );
  INVX1 U11311 ( .A(n8424), .Y(n8916) );
  INVX1 U11312 ( .A(n8425), .Y(n8917) );
  BUFX2 U11313 ( .A(n9059), .Y(n9273) );
  BUFX2 U11314 ( .A(n9059), .Y(n9272) );
  BUFX2 U11315 ( .A(n9059), .Y(n9271) );
  BUFX2 U11316 ( .A(n9058), .Y(n9270) );
  BUFX2 U11317 ( .A(n9058), .Y(n9269) );
  BUFX2 U11318 ( .A(n9058), .Y(n9268) );
  BUFX2 U11319 ( .A(n9057), .Y(n9267) );
  BUFX2 U11320 ( .A(n9057), .Y(n9266) );
  BUFX2 U11321 ( .A(n9057), .Y(n9265) );
  BUFX2 U11322 ( .A(n9056), .Y(n9264) );
  BUFX2 U11323 ( .A(n9056), .Y(n9263) );
  BUFX2 U11324 ( .A(n9056), .Y(n9262) );
  BUFX2 U11325 ( .A(n9055), .Y(n9261) );
  BUFX2 U11326 ( .A(n9055), .Y(n9260) );
  BUFX2 U11327 ( .A(n9055), .Y(n9259) );
  BUFX2 U11328 ( .A(n9054), .Y(n9258) );
  BUFX2 U11329 ( .A(n9054), .Y(n9257) );
  BUFX2 U11330 ( .A(n9054), .Y(n9256) );
  BUFX2 U11331 ( .A(n9053), .Y(n9255) );
  BUFX2 U11332 ( .A(n9053), .Y(n9254) );
  BUFX2 U11333 ( .A(n9053), .Y(n9253) );
  BUFX2 U11334 ( .A(n9052), .Y(n9252) );
  BUFX2 U11335 ( .A(n9052), .Y(n9251) );
  BUFX2 U11336 ( .A(n9052), .Y(n9250) );
  BUFX2 U11337 ( .A(n9051), .Y(n9249) );
  BUFX2 U11338 ( .A(n9051), .Y(n9248) );
  BUFX2 U11339 ( .A(n9051), .Y(n9247) );
  BUFX2 U11340 ( .A(n9050), .Y(n9246) );
  BUFX2 U11341 ( .A(n9050), .Y(n9245) );
  BUFX2 U11342 ( .A(n9050), .Y(n9244) );
  BUFX2 U11343 ( .A(n9049), .Y(n9243) );
  BUFX2 U11344 ( .A(n9049), .Y(n9242) );
  BUFX2 U11345 ( .A(n9049), .Y(n9241) );
  BUFX2 U11346 ( .A(n9048), .Y(n9240) );
  BUFX2 U11347 ( .A(n9048), .Y(n9239) );
  BUFX2 U11348 ( .A(n9048), .Y(n9238) );
  BUFX2 U11349 ( .A(n9047), .Y(n9237) );
  BUFX2 U11350 ( .A(n9047), .Y(n9236) );
  BUFX2 U11351 ( .A(n9047), .Y(n9235) );
  BUFX2 U11352 ( .A(n9046), .Y(n9234) );
  BUFX2 U11353 ( .A(n9046), .Y(n9233) );
  BUFX2 U11354 ( .A(n9046), .Y(n9232) );
  BUFX2 U11355 ( .A(n9045), .Y(n9231) );
  BUFX2 U11356 ( .A(n9045), .Y(n9230) );
  BUFX2 U11357 ( .A(n9045), .Y(n9229) );
  BUFX2 U11358 ( .A(n9044), .Y(n9228) );
  BUFX2 U11359 ( .A(n9044), .Y(n9227) );
  BUFX2 U11360 ( .A(n9044), .Y(n9226) );
  BUFX2 U11361 ( .A(n9043), .Y(n9225) );
  BUFX2 U11362 ( .A(n9043), .Y(n9224) );
  BUFX2 U11363 ( .A(n9043), .Y(n9223) );
  AND2X1 U11364 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n825 ), 
        .B(n8880), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n860 )
         );
  INVX1 U11365 ( .A(n8922), .Y(n8921) );
  INVX1 U11366 ( .A(n8920), .Y(n8919) );
  INVX1 U11367 ( .A(n8998), .Y(n8982) );
  INVX1 U11368 ( .A(n8998), .Y(n8983) );
  INVX1 U11369 ( .A(n8998), .Y(n8984) );
  INVX1 U11370 ( .A(n8998), .Y(n8985) );
  INVX1 U11371 ( .A(n9000), .Y(n8986) );
  INVX1 U11372 ( .A(n8998), .Y(n8989) );
  INVX1 U11373 ( .A(n9005), .Y(n8988) );
  INVX1 U11374 ( .A(n8998), .Y(n8987) );
  AND2X1 U11375 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .B(n9813), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n377 )
         );
  INVX1 U11376 ( .A(n8998), .Y(n8981) );
  INVX1 U11377 ( .A(p_1_cast_fu_1031_p1_31), .Y(n9490) );
  INVX1 U11378 ( .A(p_cast_fu_688_p1_31), .Y(n9540) );
  INVX1 U11379 ( .A(n8959), .Y(n8954) );
  INVX1 U11380 ( .A(n8959), .Y(n8953) );
  INVX1 U11381 ( .A(n8968), .Y(n8966) );
  INVX1 U11382 ( .A(n8968), .Y(n8965) );
  INVX1 U11383 ( .A(n9013), .Y(n9012) );
  INVX1 U11384 ( .A(n8658), .Y(n8968) );
  INVX1 U11385 ( .A(n8658), .Y(n8969) );
  INVX1 U11386 ( .A(n8658), .Y(n8970) );
  INVX1 U11387 ( .A(n8655), .Y(n8956) );
  INVX1 U11388 ( .A(n8655), .Y(n8957) );
  INVX1 U11389 ( .A(n8655), .Y(n8958) );
  INVX1 U11390 ( .A(n8655), .Y(n8959) );
  INVX1 U11391 ( .A(n8655), .Y(n8960) );
  INVX1 U11392 ( .A(n9014), .Y(n9039) );
  INVX1 U11393 ( .A(n9014), .Y(n9038) );
  INVX1 U11394 ( .A(n9014), .Y(n9037) );
  INVX1 U11395 ( .A(n9020), .Y(n9015) );
  INVX1 U11396 ( .A(n9020), .Y(n9016) );
  INVX1 U11397 ( .A(n9020), .Y(n9017) );
  INVX1 U11398 ( .A(n8956), .Y(n8955) );
  INVX1 U11399 ( .A(n9020), .Y(n9018) );
  INVX1 U11400 ( .A(n9020), .Y(n9019) );
  AND2X1 U11401 ( .A(ap_CS_fsm[12]), .B(ap_rst_n), .Y(N111) );
  AND2X1 U11402 ( .A(n970), .B(ap_rst_n), .Y(N108) );
  AND2X1 U11403 ( .A(ap_CS_fsm[7]), .B(ap_rst_n), .Y(N106) );
  AND2X1 U11404 ( .A(n1646), .B(ap_rst_n), .Y(N103) );
  AND2X1 U11405 ( .A(n8967), .B(ap_rst_n), .Y(N99) );
  INVX1 U11406 ( .A(n8970), .Y(n8967) );
  AND2X1 U11407 ( .A(\Decision_AXILiteS_s_axi_U/n247 ), .B(
        \Decision_AXILiteS_s_axi_U/n248 ), .Y(\Decision_AXILiteS_s_axi_U/n211 ) );
  BUFX2 U11408 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n14 ), 
        .Y(n8880) );
  AND2X1 U11409 ( .A(\Decision_AXILiteS_s_axi_U/n473 ), .B(
        \Decision_AXILiteS_s_axi_U/n565 ), .Y(\Decision_AXILiteS_s_axi_U/n471 ) );
  AND2X1 U11410 ( .A(n8882), .B(\Decision_AXILiteS_s_axi_U/n565 ), .Y(
        \Decision_AXILiteS_s_axi_U/n513 ) );
  AND2X1 U11411 ( .A(n8881), .B(\Decision_AXILiteS_s_axi_U/n565 ), .Y(
        \Decision_AXILiteS_s_axi_U/n408 ) );
  AND2X1 U11412 ( .A(\Decision_AXILiteS_s_axi_U/n351 ), .B(
        \Decision_AXILiteS_s_axi_U/n565 ), .Y(\Decision_AXILiteS_s_axi_U/n354 ) );
  INVX1 U11413 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n370 ), 
        .Y(n9815) );
  INVX1 U11414 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n375 ), 
        .Y(n9818) );
  INVX1 U11415 ( .A(n8405), .Y(n10276) );
  INVX1 U11416 ( .A(n8396), .Y(n9994) );
  OR2X1 U11417 ( .A(N472), .B(ap_CS_fsm[1]), .Y(n8423) );
  INVX1 U11418 ( .A(n8423), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n7 ) );
  INVX1 U11419 ( .A(n11793), .Y(n9345) );
  INVX1 U11420 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n410 ), 
        .Y(n9813) );
  BUFX2 U11421 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n17 ), 
        .Y(n8877) );
  INVX1 U11422 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n372 ), 
        .Y(n9817) );
  BUFX2 U11423 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n17 ), 
        .Y(n8876) );
  BUFX2 U11424 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n37 ), .Y(n8870) );
  BUFX2 U11425 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n35 ), .Y(n8873) );
  INVX1 U11426 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n671 ), 
        .Y(n8904) );
  INVX1 U11427 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n652 ), 
        .Y(n8902) );
  INVX1 U11428 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n740 ), 
        .Y(n8912) );
  INVX1 U11429 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n723 ), 
        .Y(n8910) );
  INVX1 U11430 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n757 ), 
        .Y(n8914) );
  AND2X1 U11431 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n825 ), 
        .B(n8878), .Y(n8424) );
  AND2X1 U11432 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n825 ), 
        .B(n8879), .Y(n8425) );
  AND2X1 U11433 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .B(n4692), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n670 )
         );
  AND2X1 U11434 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n352 ), 
        .B(n9809), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n688 )
         );
  AND2X1 U11435 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n354 ), 
        .B(n9809), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n669 )
         );
  INVX1 U11436 ( .A(n8100), .Y(n9993) );
  AND2X1 U11437 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n352 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 ), .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n32 ) );
  AND2X1 U11438 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n354 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n360 ), .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n31 ) );
  INVX1 U11439 ( .A(n8908), .Y(n8907) );
  INVX1 U11440 ( .A(n8906), .Y(n8905) );
  INVX1 U11441 ( .A(n8900), .Y(n8899) );
  AND2X1 U11442 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n352 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 ), .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n25 ) );
  AND2X1 U11443 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n354 ), 
        .B(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n353 ), .Y(\recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n24 ) );
  AND2X1 U11444 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n670 ), 
        .B(n4693), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n825 )
         );
  INVX1 U11445 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n650 ), 
        .Y(n9470) );
  INVX1 U11446 ( .A(n7631), .Y(n10896) );
  INVX1 U11447 ( .A(p_1_cast_fu_1031_p1[1]), .Y(n9480) );
  INVX1 U11448 ( .A(p_cast_fu_688_p1[1]), .Y(n9536) );
  INVX1 U11449 ( .A(n11511), .Y(n9749) );
  INVX1 U11450 ( .A(n11769), .Y(n9330) );
  INVX1 U11451 ( .A(n1230), .Y(n10243) );
  INVX1 U11452 ( .A(n1800), .Y(n9935) );
  INVX1 U11453 ( .A(n11694), .Y(n9641) );
  INVX1 U11454 ( .A(n12158), .Y(n9760) );
  INVX1 U11455 ( .A(n11680), .Y(n9628) );
  INVX1 U11456 ( .A(n12144), .Y(n9745) );
  INVX1 U11457 ( .A(n11535), .Y(n9715) );
  INVX1 U11458 ( .A(n11704), .Y(n9600) );
  INVX1 U11459 ( .A(n12168), .Y(n9711) );
  INVX1 U11460 ( .A(n8063), .Y(n9692) );
  INVX1 U11461 ( .A(CircularBuffer_len_read_assign_3_fu_1091_p3[3]), .Y(n10537) );
  INVX1 U11462 ( .A(CircularBuffer_len_read_assign_1_fu_778_p3[3]), .Y(n10072)
         );
  BUFX2 U11463 ( .A(n9061), .Y(n9059) );
  BUFX2 U11464 ( .A(n9061), .Y(n9058) );
  BUFX2 U11465 ( .A(n9062), .Y(n9057) );
  BUFX2 U11466 ( .A(n9062), .Y(n9056) );
  BUFX2 U11467 ( .A(n9062), .Y(n9055) );
  BUFX2 U11468 ( .A(n9063), .Y(n9054) );
  BUFX2 U11469 ( .A(n9063), .Y(n9053) );
  BUFX2 U11470 ( .A(n9063), .Y(n9052) );
  BUFX2 U11471 ( .A(n9064), .Y(n9051) );
  BUFX2 U11472 ( .A(n9064), .Y(n9050) );
  BUFX2 U11473 ( .A(n9064), .Y(n9049) );
  BUFX2 U11474 ( .A(n9065), .Y(n9048) );
  BUFX2 U11475 ( .A(n9065), .Y(n9047) );
  BUFX2 U11476 ( .A(n9065), .Y(n9046) );
  BUFX2 U11477 ( .A(n9066), .Y(n9045) );
  BUFX2 U11478 ( .A(n9066), .Y(n9044) );
  BUFX2 U11479 ( .A(n9066), .Y(n9043) );
  BUFX2 U11480 ( .A(n9060), .Y(n9274) );
  BUFX2 U11481 ( .A(n9061), .Y(n9060) );
  INVX1 U11482 ( .A(n8428), .Y(n8972) );
  AND2X1 U11483 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .B(n9811), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n446 )
         );
  AND2X1 U11484 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .B(n9812), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n412 )
         );
  AND2X1 U11485 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n44 ), 
        .B(n9810), .Y(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n480 )
         );
  INVX1 U11486 ( .A(n8998), .Y(n8997) );
  INVX1 U11487 ( .A(n8998), .Y(n8996) );
  INVX1 U11488 ( .A(n9001), .Y(n8995) );
  INVX1 U11489 ( .A(n9003), .Y(n8994) );
  INVX1 U11490 ( .A(n8998), .Y(n8992) );
  INVX1 U11491 ( .A(n9002), .Y(n8993) );
  INVX1 U11492 ( .A(ap_CS_fsm[1]), .Y(n8978) );
  INVX1 U11493 ( .A(n8999), .Y(n8990) );
  INVX1 U11494 ( .A(ap_CS_fsm[1]), .Y(n8977) );
  INVX1 U11495 ( .A(n8429), .Y(n8883) );
  INVX1 U11496 ( .A(n3149), .Y(n8922) );
  INVX1 U11497 ( .A(n3151), .Y(n8920) );
  INVX1 U11498 ( .A(n8998), .Y(n8991) );
  INVX1 U11499 ( .A(CircularBuffer_len_read_assign_3_fu_1091_p3[1]), .Y(n10539) );
  INVX1 U11500 ( .A(CircularBuffer_len_read_assign_1_fu_778_p3[1]), .Y(n10074)
         );
  INVX1 U11501 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n615 ), 
        .Y(n9468) );
  INVX1 U11502 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n547 ), 
        .Y(n9467) );
  INVX1 U11503 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n807 ), 
        .Y(n9466) );
  INVX1 U11504 ( .A(ap_CS_fsm[4]), .Y(n8998) );
  INVX1 U11505 ( .A(ap_CS_fsm[4]), .Y(n8999) );
  INVX1 U11506 ( .A(ap_CS_fsm[4]), .Y(n9000) );
  INVX1 U11507 ( .A(ap_CS_fsm[4]), .Y(n9001) );
  INVX1 U11508 ( .A(ap_CS_fsm[4]), .Y(n9002) );
  INVX1 U11509 ( .A(ap_CS_fsm[4]), .Y(n9003) );
  INVX1 U11510 ( .A(ap_CS_fsm[4]), .Y(n9004) );
  AND2X1 U11511 ( .A(n9310), .B(\Decision_AXILiteS_s_axi_U/n248 ), .Y(
        \Decision_AXILiteS_s_axi_U/n159 ) );
  INVX1 U11512 ( .A(ap_CS_fsm[4]), .Y(n9005) );
  INVX1 U11513 ( .A(ap_CS_fsm[4]), .Y(n9006) );
  INVX1 U11514 ( .A(ap_CS_fsm[4]), .Y(n9008) );
  INVX1 U11515 ( .A(ap_CS_fsm[4]), .Y(n9009) );
  INVX1 U11516 ( .A(ap_CS_fsm[4]), .Y(n9010) );
  INVX1 U11517 ( .A(ap_CS_fsm[4]), .Y(n9007) );
  INVX1 U11518 ( .A(CircularBuffer_len_read_assign_3_fu_1091_p3[2]), .Y(n10538) );
  INVX1 U11519 ( .A(CircularBuffer_len_read_assign_1_fu_778_p3[2]), .Y(n10073)
         );
  AND2X1 U11520 ( .A(\Decision_AXILiteS_s_axi_U/n248 ), .B(n9309), .Y(
        \Decision_AXILiteS_s_axi_U/n158 ) );
  INVX1 U11521 ( .A(CircularBuffer_len_read_assign_3_fu_1091_p3[4]), .Y(n10536) );
  INVX1 U11522 ( .A(CircularBuffer_len_read_assign_1_fu_778_p3[4]), .Y(n10071)
         );
  INVX1 U11523 ( .A(ap_CS_fsm[13]), .Y(n8896) );
  INVX1 U11524 ( .A(n2872), .Y(n8923) );
  INVX1 U11525 ( .A(ap_CS_fsm[7]), .Y(n9013) );
  INVX1 U11526 ( .A(n9020), .Y(n9014) );
  INVX1 U11527 ( .A(n8658), .Y(n8971) );
  INVX1 U11528 ( .A(ap_CS_fsm[12]), .Y(n9041) );
  AND2X1 U11529 ( .A(n8976), .B(ap_rst_n), .Y(N100) );
  INVX1 U11530 ( .A(i_8_fu_1148_p2[31]), .Y(n10306) );
  INVX1 U11531 ( .A(i_2_fu_823_p2[31]), .Y(n9965) );
  INVX1 U11532 ( .A(n2200), .Y(n9995) );
  INVX1 U11533 ( .A(i_5_fu_854_p2[1]), .Y(n10023) );
  INVX1 U11534 ( .A(n2194), .Y(n10277) );
  INVX1 U11535 ( .A(i_11_fu_1179_p2[1]), .Y(n10305) );
  BUFX2 U11536 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n13 ), 
        .Y(n8879) );
  INVX1 U11537 ( .A(n11780), .Y(n9324) );
  INVX1 U11538 ( .A(n11522), .Y(n9764) );
  INVX1 U11539 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n479 ), 
        .Y(n9811) );
  AND2X1 U11540 ( .A(n9318), .B(\Decision_AXILiteS_s_axi_U/n248 ), .Y(
        \Decision_AXILiteS_s_axi_U/n210 ) );
  AND2X1 U11541 ( .A(n9011), .B(n10056), .Y(n373) );
  AND2X1 U11542 ( .A(n10534), .B(n9040), .Y(n387) );
  AND2X1 U11543 ( .A(\Decision_AXILiteS_s_axi_U/n533 ), .B(
        \Decision_AXILiteS_s_axi_U/n565 ), .Y(\Decision_AXILiteS_s_axi_U/n555 ) );
  AND2X1 U11544 ( .A(\Decision_AXILiteS_s_axi_U/n429 ), .B(
        \Decision_AXILiteS_s_axi_U/n565 ), .Y(\Decision_AXILiteS_s_axi_U/n450 ) );
  OR2X1 U11545 ( .A(n9638), .B(sum_1_phi_fu_379_p4[28]), .Y(n11767) );
  OR2X1 U11546 ( .A(n9755), .B(sum_phi_fu_311_p4[28]), .Y(n11509) );
  OR2X1 U11547 ( .A(n9636), .B(n2245), .Y(n11678) );
  OR2X1 U11548 ( .A(n9753), .B(n2738), .Y(n12142) );
  OR2X1 U11549 ( .A(p_tmp_i_fu_587_p3[3]), .B(p_tmp_i_fu_587_p3[5]), .Y(n1947)
         );
  INVX1 U11550 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n373 ), 
        .Y(n9819) );
  INVX1 U11551 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n363 ), 
        .Y(n9820) );
  INVX1 U11552 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n445 ), 
        .Y(n9812) );
  INVX1 U11553 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n513 ), 
        .Y(n9810) );
  OR2X1 U11554 ( .A(n9773), .B(p_1_cast_fu_1031_p1[12]), .Y(n11582) );
  OR2X1 U11555 ( .A(n9512), .B(p_cast_fu_688_p1[12]), .Y(n12215) );
  OR2X1 U11556 ( .A(n9586), .B(sum_1_phi_fu_379_p4[12]), .Y(n11722) );
  OR2X1 U11557 ( .A(n9693), .B(sum_phi_fu_311_p4[12]), .Y(n11464) );
  OR2X1 U11558 ( .A(n9584), .B(n2277), .Y(n11633) );
  OR2X1 U11559 ( .A(n9690), .B(n2770), .Y(n12097) );
  BUFX2 U11560 ( .A(n7252), .Y(n8885) );
  BUFX2 U11561 ( .A(n7428), .Y(n8887) );
  INVX1 U11562 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n371 ), 
        .Y(n9816) );
  INVX1 U11563 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n365 ), 
        .Y(n9814) );
  BUFX2 U11564 ( .A(n7252), .Y(n8884) );
  BUFX2 U11565 ( .A(n7428), .Y(n8886) );
  INVX1 U11566 ( .A(n11650), .Y(n9568) );
  INVX1 U11567 ( .A(n12114), .Y(n9672) );
  INVX1 U11568 ( .A(n11481), .Y(n9675) );
  AND2X1 U11569 ( .A(n11753), .B(n9560), .Y(n11754) );
  AND2X1 U11570 ( .A(n11539), .B(n9724), .Y(n11540) );
  AND2X1 U11571 ( .A(n11708), .B(n9610), .Y(n11709) );
  AND2X1 U11572 ( .A(n12172), .B(n9721), .Y(n12173) );
  BUFX2 U11573 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n15 ), 
        .Y(n8878) );
  INVX1 U11574 ( .A(\Decision_AXILiteS_s_axi_U/n320 ), .Y(n9315) );
  INVX1 U11575 ( .A(n11580), .Y(n9484) );
  INVX1 U11576 ( .A(n12213), .Y(n9503) );
  INVX1 U11577 ( .A(i_11_fu_1179_p2[31]), .Y(n10279) );
  INVX1 U11578 ( .A(i_5_fu_854_p2[31]), .Y(n9997) );
  INVX1 U11579 ( .A(\Decision_AXILiteS_s_axi_U/n322 ), .Y(n9314) );
  INVX1 U11580 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n15 ), .Y(n10275) );
  INVX1 U11581 ( .A(n5971), .Y(n9809) );
  BUFX2 U11582 ( .A(\Decision_AXILiteS_s_axi_U/n492 ), .Y(n8882) );
  BUFX2 U11583 ( .A(\Decision_AXILiteS_s_axi_U/n383 ), .Y(n8881) );
  INVX1 U11584 ( .A(\dp_cluster_0/N954 ), .Y(n10776) );
  INVX1 U11585 ( .A(\dp_cluster_1/N922 ), .Y(n10742) );
  OR2X1 U11586 ( .A(\Decision_AXILiteS_s_axi_U/n315 ), .B(n8918), .Y(n8426) );
  INVX1 U11587 ( .A(n8426), .Y(\Decision_AXILiteS_s_axi_U/n248 ) );
  INVX1 U11588 ( .A(n11882), .Y(n10413) );
  INVX1 U11589 ( .A(n11158), .Y(n10497) );
  INVX1 U11590 ( .A(n12079), .Y(n9709) );
  INVX1 U11591 ( .A(n11990), .Y(n9602) );
  OR2X1 U11592 ( .A(n9598), .B(sum_1_phi_fu_379_p4[16]), .Y(n11763) );
  INVX1 U11593 ( .A(n11739), .Y(n9352) );
  INVX1 U11594 ( .A(n11894), .Y(n10430) );
  INVX1 U11595 ( .A(n11170), .Y(n10514) );
  INVX1 U11596 ( .A(n12091), .Y(n9736) );
  INVX1 U11597 ( .A(n12002), .Y(n9623) );
  INVX1 U11598 ( .A(n11805), .Y(n9322) );
  INVX1 U11599 ( .A(n11567), .Y(n9481) );
  INVX1 U11600 ( .A(n12200), .Y(n9498) );
  INVX1 U11601 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n361 ), 
        .Y(n9821) );
  INVX1 U11602 ( .A(n11726), .Y(n9366) );
  INVX1 U11603 ( .A(n11729), .Y(n9362) );
  INVX1 U11604 ( .A(n11776), .Y(n9331) );
  INVX1 U11605 ( .A(n11468), .Y(n9676) );
  INVX1 U11606 ( .A(n11471), .Y(n9686) );
  INVX1 U11607 ( .A(n11518), .Y(n9750) );
  INVX1 U11608 ( .A(n11687), .Y(n9629) );
  INVX1 U11609 ( .A(n12151), .Y(n9746) );
  INVX1 U11610 ( .A(n11637), .Y(n9569) );
  INVX1 U11611 ( .A(n11640), .Y(n9576) );
  INVX1 U11612 ( .A(n12101), .Y(n9673) );
  INVX1 U11613 ( .A(n12104), .Y(n9682) );
  INVX1 U11614 ( .A(n11586), .Y(n9486) );
  INVX1 U11615 ( .A(n11589), .Y(n9474) );
  INVX1 U11616 ( .A(n11596), .Y(n9478) );
  INVX1 U11617 ( .A(n12219), .Y(n9506) );
  INVX1 U11618 ( .A(n12222), .Y(n9509) );
  INVX1 U11619 ( .A(n12229), .Y(n9515) );
  BUFX2 U11620 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n55 ), .Y(n8871) );
  BUFX2 U11621 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n53 ), .Y(n8874) );
  BUFX2 U11622 ( .A(\recentVBools_data_U/Decision_recentVBools_data_ram_U/n64 ), .Y(n8875) );
  BUFX2 U11623 ( .A(\recentABools_data_U/Decision_recentVBools_data_ram_U/n66 ), .Y(n8872) );
  INVX1 U11624 ( .A(n8858), .Y(n9320) );
  INVX1 U11625 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n706 ), 
        .Y(n8908) );
  INVX1 U11626 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n689 ), 
        .Y(n8906) );
  INVX1 U11627 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n550 ), 
        .Y(n8900) );
  INVX1 U11628 ( .A(n11716), .Y(n9622) );
  INVX1 U11629 ( .A(n12180), .Y(n9737) );
  INVX1 U11630 ( .A(n11547), .Y(n9740) );
  INVX1 U11631 ( .A(\Decision_AXILiteS_s_axi_U/n631 ), .Y(n9316) );
  INVX1 U11632 ( .A(n8427), .Y(\Decision_AXILiteS_s_axi_U/n351 ) );
  INVX1 U11633 ( .A(\Decision_AXILiteS_s_axi_U/n340 ), .Y(n9309) );
  INVX1 U11634 ( .A(\Decision_AXILiteS_s_axi_U/n339 ), .Y(n9310) );
  INVX1 U11635 ( .A(n8978), .Y(n8976) );
  INVX1 U11636 ( .A(n8978), .Y(n8975) );
  INVX1 U11637 ( .A(n7434), .Y(n9279) );
  AND2X1 U11638 ( .A(n9319), .B(n9317), .Y(\Decision_AXILiteS_s_axi_U/n310 )
         );
  INVX1 U11639 ( .A(n365), .Y(n9824) );
  OR2X1 U11640 ( .A(n8922), .B(CircularBuffer_len_read_assign_2_fu_1085_p2[2]), 
        .Y(CircularBuffer_len_read_assign_3_fu_1091_p3[2]) );
  OR2X1 U11641 ( .A(n8920), .B(CircularBuffer_len_read_assign_fu_772_p2[2]), 
        .Y(CircularBuffer_len_read_assign_1_fu_778_p3[2]) );
  OR2X1 U11642 ( .A(n8922), .B(CircularBuffer_len_read_assign_2_fu_1085_p2[4]), 
        .Y(CircularBuffer_len_read_assign_3_fu_1091_p3[4]) );
  OR2X1 U11643 ( .A(n8920), .B(CircularBuffer_len_read_assign_fu_772_p2[4]), 
        .Y(CircularBuffer_len_read_assign_1_fu_778_p3[4]) );
  INVX1 U11644 ( .A(n8383), .Y(n9311) );
  INVX1 U11645 ( .A(n8888), .Y(n9823) );
  INVX1 U11646 ( .A(n5962), .Y(n9278) );
  INVX1 U11647 ( .A(i_8_fu_1148_p2[1]), .Y(n10332) );
  INVX1 U11648 ( .A(i_2_fu_823_p2[1]), .Y(n9991) );
  BUFX2 U11649 ( .A(n2050), .Y(n8869) );
  BUFX2 U11650 ( .A(n2050), .Y(n8868) );
  INVX1 U11651 ( .A(n2192), .Y(n10274) );
  INVX1 U11652 ( .A(sum_1_phi_fu_379_p4[8]), .Y(n9368) );
  INVX1 U11653 ( .A(sum_phi_fu_311_p4[8]), .Y(n10064) );
  INVX1 U11654 ( .A(n8889), .Y(n9822) );
  INVX1 U11655 ( .A(n8653), .Y(n8974) );
  INVX1 U11656 ( .A(n8654), .Y(n8973) );
  INVX1 U11657 ( .A(sum_1_phi_fu_379_p4[7]), .Y(n9371) );
  INVX1 U11658 ( .A(sum_1_phi_fu_379_p4[3]), .Y(n9377) );
  INVX1 U11659 ( .A(sum_1_phi_fu_379_p4[11]), .Y(n9363) );
  INVX1 U11660 ( .A(sum_1_phi_fu_379_p4[15]), .Y(n9356) );
  INVX1 U11661 ( .A(sum_phi_fu_311_p4[11]), .Y(n10065) );
  INVX1 U11662 ( .A(sum_phi_fu_311_p4[15]), .Y(n10066) );
  INVX1 U11663 ( .A(sum_phi_fu_311_p4[23]), .Y(n10068) );
  INVX1 U11664 ( .A(sum_1_phi_fu_379_p4[19]), .Y(n9347) );
  INVX1 U11665 ( .A(sum_phi_fu_311_p4[7]), .Y(n10063) );
  INVX1 U11666 ( .A(sum_phi_fu_311_p4[27]), .Y(n10069) );
  INVX1 U11667 ( .A(sum_phi_fu_311_p4[19]), .Y(n10067) );
  INVX1 U11668 ( .A(sum_1_phi_fu_379_p4[27]), .Y(n9332) );
  INVX1 U11669 ( .A(sum_phi_fu_311_p4[3]), .Y(n10062) );
  INVX1 U11670 ( .A(sum_1_phi_fu_379_p4[23]), .Y(n9340) );
  INVX1 U11671 ( .A(n12055), .Y(n9743) );
  INVX1 U11672 ( .A(n11966), .Y(n9630) );
  INVX1 U11673 ( .A(n12069), .Y(n9758) );
  INVX1 U11674 ( .A(n11980), .Y(n9643) );
  INVX1 U11675 ( .A(n11736), .Y(n9355) );
  INVX1 U11676 ( .A(n11478), .Y(n9702) );
  INVX1 U11677 ( .A(n11825), .Y(n10404) );
  INVX1 U11678 ( .A(n11647), .Y(n9589) );
  INVX1 U11679 ( .A(n12111), .Y(n9698) );
  INVX1 U11680 ( .A(n12022), .Y(n9696) );
  INVX1 U11681 ( .A(n11933), .Y(n9591) );
  INVX1 U11682 ( .A(n11872), .Y(n10446) );
  INVX1 U11683 ( .A(n11148), .Y(n10530) );
  INVX1 U11684 ( .A(n11858), .Y(n10435) );
  INVX1 U11685 ( .A(n11134), .Y(n10519) );
  INVX1 U11686 ( .A(n11101), .Y(n10488) );
  OR2X1 U11687 ( .A(n8922), .B(CircularBuffer_len_read_assign_2_fu_1085_p2[1]), 
        .Y(CircularBuffer_len_read_assign_3_fu_1091_p3[1]) );
  OR2X1 U11688 ( .A(n8920), .B(CircularBuffer_len_read_assign_fu_772_p2[1]), 
        .Y(CircularBuffer_len_read_assign_1_fu_778_p3[1]) );
  INVX1 U11689 ( .A(p_1_cast_fu_1031_p1[8]), .Y(n9487) );
  INVX1 U11690 ( .A(p_cast_fu_688_p1[8]), .Y(n9539) );
  INVX1 U11691 ( .A(n8657), .Y(n8930) );
  INVX1 U11692 ( .A(n8656), .Y(n8929) );
  OR2X1 U11693 ( .A(n9592), .B(sum_1_phi_fu_379_p4[13]), .Y(n11732) );
  OR2X1 U11694 ( .A(n9699), .B(sum_phi_fu_311_p4[13]), .Y(n11474) );
  OR2X1 U11695 ( .A(n9761), .B(sum_phi_fu_311_p4[29]), .Y(n11521) );
  OR2X1 U11696 ( .A(n9644), .B(sum_1_phi_fu_379_p4[29]), .Y(n11779) );
  INVX1 U11697 ( .A(n11617), .Y(n9489) );
  INVX1 U11698 ( .A(n12250), .Y(n9532) );
  XNOR2X1 U11699 ( .A(n8665), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[1]), 
        .Y(n8430) );
  XNOR2X1 U11700 ( .A(n8504), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[2]), 
        .Y(n8431) );
  XNOR2X1 U11701 ( .A(n8506), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[3]), 
        .Y(n8432) );
  XNOR2X1 U11702 ( .A(n8508), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[4]), 
        .Y(n8433) );
  XNOR2X1 U11703 ( .A(n8510), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[5]), 
        .Y(n8434) );
  XNOR2X1 U11704 ( .A(n8512), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[6]), 
        .Y(n8435) );
  XNOR2X1 U11705 ( .A(n8514), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[7]), 
        .Y(n8436) );
  XNOR2X1 U11706 ( .A(n8516), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[8]), 
        .Y(n8437) );
  XNOR2X1 U11707 ( .A(n8518), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[9]), 
        .Y(n8438) );
  XNOR2X1 U11708 ( .A(n8520), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[10]), 
        .Y(n8439) );
  XNOR2X1 U11709 ( .A(n8490), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[11]), 
        .Y(n8440) );
  XNOR2X1 U11710 ( .A(n8522), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[12]), 
        .Y(n8441) );
  XNOR2X1 U11711 ( .A(n8492), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[13]), 
        .Y(n8442) );
  XNOR2X1 U11712 ( .A(n8494), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[14]), 
        .Y(n8443) );
  XNOR2X1 U11713 ( .A(n8496), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[15]), 
        .Y(n8444) );
  XNOR2X1 U11714 ( .A(n8498), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[16]), 
        .Y(n8445) );
  XNOR2X1 U11715 ( .A(n8500), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[17]), 
        .Y(n8446) );
  XNOR2X1 U11716 ( .A(n8502), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[18]), 
        .Y(n8447) );
  XNOR2X1 U11717 ( .A(n8524), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[19]), 
        .Y(n8448) );
  XNOR2X1 U11718 ( .A(n8526), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[20]), 
        .Y(n8449) );
  XNOR2X1 U11719 ( .A(n8528), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[21]), 
        .Y(n8450) );
  XNOR2X1 U11720 ( .A(n8530), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[22]), 
        .Y(n8451) );
  XNOR2X1 U11721 ( .A(n8532), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[23]), 
        .Y(n8452) );
  XNOR2X1 U11722 ( .A(n8534), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[24]), 
        .Y(n8453) );
  XNOR2X1 U11723 ( .A(n8536), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[25]), 
        .Y(n8454) );
  XNOR2X1 U11724 ( .A(n8538), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[26]), 
        .Y(n8455) );
  XNOR2X1 U11725 ( .A(n8540), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[27]), 
        .Y(n8456) );
  XNOR2X1 U11726 ( .A(n8542), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[28]), 
        .Y(n8457) );
  XNOR2X1 U11727 ( .A(n8544), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[29]), 
        .Y(n8458) );
  XNOR2X1 U11728 ( .A(n8547), .B(CircularBuffer_int_30_sum_i_fu_758_p3[30]), 
        .Y(n8459) );
  XNOR2X1 U11729 ( .A(n8545), .B(CircularBuffer_int_30_sum_i_fu_758_p3[29]), 
        .Y(n8460) );
  XNOR2X1 U11730 ( .A(n8543), .B(CircularBuffer_int_30_sum_i_fu_758_p3[28]), 
        .Y(n8461) );
  XNOR2X1 U11731 ( .A(n8541), .B(CircularBuffer_int_30_sum_i_fu_758_p3[27]), 
        .Y(n8462) );
  XNOR2X1 U11732 ( .A(n8539), .B(CircularBuffer_int_30_sum_i_fu_758_p3[26]), 
        .Y(n8463) );
  XNOR2X1 U11733 ( .A(n8537), .B(CircularBuffer_int_30_sum_i_fu_758_p3[25]), 
        .Y(n8464) );
  XNOR2X1 U11734 ( .A(n8535), .B(CircularBuffer_int_30_sum_i_fu_758_p3[24]), 
        .Y(n8465) );
  XNOR2X1 U11735 ( .A(n8533), .B(CircularBuffer_int_30_sum_i_fu_758_p3[23]), 
        .Y(n8466) );
  XNOR2X1 U11736 ( .A(n8531), .B(CircularBuffer_int_30_sum_i_fu_758_p3[22]), 
        .Y(n8467) );
  XNOR2X1 U11737 ( .A(n8529), .B(CircularBuffer_int_30_sum_i_fu_758_p3[21]), 
        .Y(n8468) );
  XNOR2X1 U11738 ( .A(n8527), .B(CircularBuffer_int_30_sum_i_fu_758_p3[20]), 
        .Y(n8469) );
  XNOR2X1 U11739 ( .A(n8525), .B(CircularBuffer_int_30_sum_i_fu_758_p3[19]), 
        .Y(n8470) );
  XNOR2X1 U11740 ( .A(n8503), .B(CircularBuffer_int_30_sum_i_fu_758_p3[18]), 
        .Y(n8471) );
  XNOR2X1 U11741 ( .A(n8501), .B(CircularBuffer_int_30_sum_i_fu_758_p3[17]), 
        .Y(n8472) );
  XNOR2X1 U11742 ( .A(n8499), .B(CircularBuffer_int_30_sum_i_fu_758_p3[16]), 
        .Y(n8473) );
  XNOR2X1 U11743 ( .A(n8497), .B(CircularBuffer_int_30_sum_i_fu_758_p3[15]), 
        .Y(n8474) );
  XNOR2X1 U11744 ( .A(n8495), .B(CircularBuffer_int_30_sum_i_fu_758_p3[14]), 
        .Y(n8475) );
  XNOR2X1 U11745 ( .A(n8493), .B(CircularBuffer_int_30_sum_i_fu_758_p3[13]), 
        .Y(n8476) );
  XNOR2X1 U11746 ( .A(n8523), .B(CircularBuffer_int_30_sum_i_fu_758_p3[12]), 
        .Y(n8477) );
  XNOR2X1 U11747 ( .A(n8491), .B(CircularBuffer_int_30_sum_i_fu_758_p3[11]), 
        .Y(n8478) );
  XNOR2X1 U11748 ( .A(n8521), .B(CircularBuffer_int_30_sum_i_fu_758_p3[10]), 
        .Y(n8479) );
  XNOR2X1 U11749 ( .A(n8519), .B(CircularBuffer_int_30_sum_i_fu_758_p3[9]), 
        .Y(n8480) );
  XNOR2X1 U11750 ( .A(n8517), .B(CircularBuffer_int_30_sum_i_fu_758_p3[8]), 
        .Y(n8481) );
  XNOR2X1 U11751 ( .A(n8515), .B(CircularBuffer_int_30_sum_i_fu_758_p3[7]), 
        .Y(n8482) );
  XNOR2X1 U11752 ( .A(n8513), .B(CircularBuffer_int_30_sum_i_fu_758_p3[6]), 
        .Y(n8483) );
  XNOR2X1 U11753 ( .A(n8511), .B(CircularBuffer_int_30_sum_i_fu_758_p3[5]), 
        .Y(n8484) );
  XNOR2X1 U11754 ( .A(n8509), .B(CircularBuffer_int_30_sum_i_fu_758_p3[4]), 
        .Y(n8485) );
  XNOR2X1 U11755 ( .A(n8507), .B(CircularBuffer_int_30_sum_i_fu_758_p3[3]), 
        .Y(n8486) );
  XNOR2X1 U11756 ( .A(n8505), .B(CircularBuffer_int_30_sum_i_fu_758_p3[2]), 
        .Y(n8487) );
  XNOR2X1 U11757 ( .A(n8666), .B(CircularBuffer_int_30_sum_i_fu_758_p3[1]), 
        .Y(n8488) );
  XNOR2X1 U11758 ( .A(n8546), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[30]), 
        .Y(n8489) );
  INVX1 U11759 ( .A(n11581), .Y(n9477) );
  INVX1 U11760 ( .A(n12214), .Y(n9514) );
  INVX1 U11761 ( .A(n11508), .Y(n9763) );
  INVX1 U11762 ( .A(n11766), .Y(n9323) );
  INVX1 U11763 ( .A(n11721), .Y(n9354) );
  INVX1 U11764 ( .A(n11463), .Y(n9701) );
  INVX1 U11765 ( .A(n11599), .Y(n9472) );
  INVX1 U11766 ( .A(n12232), .Y(n9505) );
  INVX1 U11767 ( .A(n11677), .Y(n9640) );
  INVX1 U11768 ( .A(n12141), .Y(n9759) );
  INVX1 U11769 ( .A(n11583), .Y(n9473) );
  INVX1 U11770 ( .A(n12216), .Y(n9508) );
  INVX1 U11771 ( .A(n11564), .Y(n9483) );
  INVX1 U11772 ( .A(n12197), .Y(n9502) );
  INVX1 U11773 ( .A(n11632), .Y(n9588) );
  INVX1 U11774 ( .A(n12096), .Y(n9697) );
  INVX1 U11775 ( .A(p_1_cast_fu_1031_p1[3]), .Y(n9482) );
  INVX1 U11776 ( .A(p_1_cast_fu_1031_p1[11]), .Y(n9475) );
  INVX1 U11777 ( .A(p_1_cast_fu_1031_p1[15]), .Y(n9479) );
  INVX1 U11778 ( .A(p_cast_fu_688_p1[3]), .Y(n9537) );
  INVX1 U11779 ( .A(p_cast_fu_688_p1[11]), .Y(n9534) );
  INVX1 U11780 ( .A(p_cast_fu_688_p1[15]), .Y(n9535) );
  INVX1 U11781 ( .A(p_1_cast_fu_1031_p1[7]), .Y(n9485) );
  INVX1 U11782 ( .A(p_cast_fu_688_p1[7]), .Y(n9538) );
  INVX1 U11783 ( .A(n11723), .Y(n9361) );
  INVX1 U11784 ( .A(n11465), .Y(n9685) );
  OR2X1 U11785 ( .A(n9604), .B(sum_1_phi_fu_379_p4[17]), .Y(n11790) );
  OR2X1 U11786 ( .A(n9618), .B(sum_1_phi_fu_379_p4[21]), .Y(n11797) );
  OR2X1 U11787 ( .A(n9730), .B(sum_phi_fu_311_p4[21]), .Y(n11539) );
  OR2X1 U11788 ( .A(n9713), .B(sum_phi_fu_311_p4[17]), .Y(n11532) );
  OR2X1 U11789 ( .A(n9747), .B(sum_phi_fu_311_p4[25]), .Y(n11514) );
  OR2X1 U11790 ( .A(n9632), .B(sum_1_phi_fu_379_p4[25]), .Y(n11772) );
  INVX1 U11791 ( .A(n11623), .Y(n9488) );
  INVX1 U11792 ( .A(n12256), .Y(n9525) );
  OR2X1 U11793 ( .A(n9774), .B(p_1_cast_fu_1031_p1[13]), .Y(n11592) );
  OR2X1 U11794 ( .A(n9513), .B(p_cast_fu_688_p1[13]), .Y(n12225) );
  BUFX2 U11795 ( .A(ap_clk), .Y(n9061) );
  BUFX2 U11796 ( .A(ap_clk), .Y(n9062) );
  BUFX2 U11797 ( .A(ap_clk), .Y(n9063) );
  BUFX2 U11798 ( .A(ap_clk), .Y(n9064) );
  BUFX2 U11799 ( .A(ap_clk), .Y(n9065) );
  BUFX2 U11800 ( .A(ap_clk), .Y(n9066) );
  INVX1 U11801 ( .A(n11634), .Y(n9575) );
  INVX1 U11802 ( .A(n12098), .Y(n9681) );
  AND2X1 U11803 ( .A(n8520), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[10]), 
        .Y(n8490) );
  AND2X1 U11804 ( .A(n8521), .B(CircularBuffer_int_30_sum_i_fu_758_p3[10]), 
        .Y(n8491) );
  AND2X1 U11805 ( .A(n8522), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[12]), 
        .Y(n8492) );
  AND2X1 U11806 ( .A(n8523), .B(CircularBuffer_int_30_sum_i_fu_758_p3[12]), 
        .Y(n8493) );
  AND2X1 U11807 ( .A(n8492), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[13]), 
        .Y(n8494) );
  AND2X1 U11808 ( .A(n8493), .B(CircularBuffer_int_30_sum_i_fu_758_p3[13]), 
        .Y(n8495) );
  AND2X1 U11809 ( .A(n8494), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[14]), 
        .Y(n8496) );
  AND2X1 U11810 ( .A(n8495), .B(CircularBuffer_int_30_sum_i_fu_758_p3[14]), 
        .Y(n8497) );
  AND2X1 U11811 ( .A(n8496), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[15]), 
        .Y(n8498) );
  AND2X1 U11812 ( .A(n8497), .B(CircularBuffer_int_30_sum_i_fu_758_p3[15]), 
        .Y(n8499) );
  AND2X1 U11813 ( .A(n8498), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[16]), 
        .Y(n8500) );
  AND2X1 U11814 ( .A(n8499), .B(CircularBuffer_int_30_sum_i_fu_758_p3[16]), 
        .Y(n8501) );
  AND2X1 U11815 ( .A(n8500), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[17]), 
        .Y(n8502) );
  AND2X1 U11816 ( .A(n8501), .B(CircularBuffer_int_30_sum_i_fu_758_p3[17]), 
        .Y(n8503) );
  AND2X1 U11817 ( .A(n8665), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[1]), 
        .Y(n8504) );
  AND2X1 U11818 ( .A(n8666), .B(CircularBuffer_int_30_sum_i_fu_758_p3[1]), .Y(
        n8505) );
  AND2X1 U11819 ( .A(n8504), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[2]), 
        .Y(n8506) );
  AND2X1 U11820 ( .A(n8505), .B(CircularBuffer_int_30_sum_i_fu_758_p3[2]), .Y(
        n8507) );
  AND2X1 U11821 ( .A(n8506), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[3]), 
        .Y(n8508) );
  AND2X1 U11822 ( .A(n8507), .B(CircularBuffer_int_30_sum_i_fu_758_p3[3]), .Y(
        n8509) );
  AND2X1 U11823 ( .A(n8508), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[4]), 
        .Y(n8510) );
  AND2X1 U11824 ( .A(n8509), .B(CircularBuffer_int_30_sum_i_fu_758_p3[4]), .Y(
        n8511) );
  AND2X1 U11825 ( .A(n8510), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[5]), 
        .Y(n8512) );
  AND2X1 U11826 ( .A(n8511), .B(CircularBuffer_int_30_sum_i_fu_758_p3[5]), .Y(
        n8513) );
  AND2X1 U11827 ( .A(n8512), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[6]), 
        .Y(n8514) );
  AND2X1 U11828 ( .A(n8513), .B(CircularBuffer_int_30_sum_i_fu_758_p3[6]), .Y(
        n8515) );
  AND2X1 U11829 ( .A(n8514), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[7]), 
        .Y(n8516) );
  AND2X1 U11830 ( .A(n8515), .B(CircularBuffer_int_30_sum_i_fu_758_p3[7]), .Y(
        n8517) );
  AND2X1 U11831 ( .A(n8516), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[8]), 
        .Y(n8518) );
  AND2X1 U11832 ( .A(n8517), .B(CircularBuffer_int_30_sum_i_fu_758_p3[8]), .Y(
        n8519) );
  AND2X1 U11833 ( .A(n8518), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[9]), 
        .Y(n8520) );
  AND2X1 U11834 ( .A(n8519), .B(CircularBuffer_int_30_sum_i_fu_758_p3[9]), .Y(
        n8521) );
  AND2X1 U11835 ( .A(n8490), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[11]), 
        .Y(n8522) );
  AND2X1 U11836 ( .A(n8491), .B(CircularBuffer_int_30_sum_i_fu_758_p3[11]), 
        .Y(n8523) );
  AND2X1 U11837 ( .A(n8502), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[18]), 
        .Y(n8524) );
  AND2X1 U11838 ( .A(n8503), .B(CircularBuffer_int_30_sum_i_fu_758_p3[18]), 
        .Y(n8525) );
  AND2X1 U11839 ( .A(n8524), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[19]), 
        .Y(n8526) );
  AND2X1 U11840 ( .A(n8525), .B(CircularBuffer_int_30_sum_i_fu_758_p3[19]), 
        .Y(n8527) );
  AND2X1 U11841 ( .A(n8526), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[20]), 
        .Y(n8528) );
  AND2X1 U11842 ( .A(n8527), .B(CircularBuffer_int_30_sum_i_fu_758_p3[20]), 
        .Y(n8529) );
  AND2X1 U11843 ( .A(n8528), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[21]), 
        .Y(n8530) );
  AND2X1 U11844 ( .A(n8529), .B(CircularBuffer_int_30_sum_i_fu_758_p3[21]), 
        .Y(n8531) );
  AND2X1 U11845 ( .A(n8530), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[22]), 
        .Y(n8532) );
  AND2X1 U11846 ( .A(n8531), .B(CircularBuffer_int_30_sum_i_fu_758_p3[22]), 
        .Y(n8533) );
  AND2X1 U11847 ( .A(n8532), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[23]), 
        .Y(n8534) );
  AND2X1 U11848 ( .A(n8533), .B(CircularBuffer_int_30_sum_i_fu_758_p3[23]), 
        .Y(n8535) );
  AND2X1 U11849 ( .A(n8534), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[24]), 
        .Y(n8536) );
  AND2X1 U11850 ( .A(n8535), .B(CircularBuffer_int_30_sum_i_fu_758_p3[24]), 
        .Y(n8537) );
  AND2X1 U11851 ( .A(n8536), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[25]), 
        .Y(n8538) );
  AND2X1 U11852 ( .A(n8537), .B(CircularBuffer_int_30_sum_i_fu_758_p3[25]), 
        .Y(n8539) );
  AND2X1 U11853 ( .A(n8538), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[26]), 
        .Y(n8540) );
  AND2X1 U11854 ( .A(n8539), .B(CircularBuffer_int_30_sum_i_fu_758_p3[26]), 
        .Y(n8541) );
  AND2X1 U11855 ( .A(n8540), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[27]), 
        .Y(n8542) );
  AND2X1 U11856 ( .A(n8541), .B(CircularBuffer_int_30_sum_i_fu_758_p3[27]), 
        .Y(n8543) );
  AND2X1 U11857 ( .A(n8542), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[28]), 
        .Y(n8544) );
  AND2X1 U11858 ( .A(n8543), .B(CircularBuffer_int_30_sum_i_fu_758_p3[28]), 
        .Y(n8545) );
  AND2X1 U11859 ( .A(n8544), .B(CircularBuffer_int_30_sum_i1_fu_1071_p3[29]), 
        .Y(n8546) );
  AND2X1 U11860 ( .A(n8545), .B(CircularBuffer_int_30_sum_i_fu_758_p3[29]), 
        .Y(n8547) );
  INVX1 U11861 ( .A(n8857), .Y(n9321) );
  OR2X1 U11862 ( .A(n9564), .B(sum_1_phi_fu_379_p4[5]), .Y(n11753) );
  OR2X1 U11863 ( .A(n9665), .B(sum_phi_fu_311_p4[5]), .Y(n11495) );
  INVX1 U11864 ( .A(n11765), .Y(n9337) );
  OR2X1 U11865 ( .A(n9612), .B(sum_1_phi_fu_379_p4[20]), .Y(n11764) );
  INVX1 U11866 ( .A(n11800), .Y(n9338) );
  INVX1 U11867 ( .A(n11507), .Y(n9723) );
  OR2X1 U11868 ( .A(n9724), .B(sum_phi_fu_311_p4[20]), .Y(n11506) );
  INVX1 U11869 ( .A(n11542), .Y(n9732) );
  AND2X1 U11870 ( .A(n473), .B(n474), .Y(n439) );
  AND2X1 U11871 ( .A(n431), .B(n432), .Y(n397) );
  INVX1 U11872 ( .A(n11676), .Y(n9608) );
  OR2X1 U11873 ( .A(n9610), .B(n2261), .Y(n11675) );
  INVX1 U11874 ( .A(n11711), .Y(n9614) );
  INVX1 U11875 ( .A(n12140), .Y(n9720) );
  OR2X1 U11876 ( .A(n9721), .B(n2754), .Y(n12139) );
  INVX1 U11877 ( .A(n12175), .Y(n9728) );
  OR2X1 U11878 ( .A(n9586), .B(n2275), .Y(n11643) );
  OR2X1 U11879 ( .A(n9693), .B(n2768), .Y(n12107) );
  OR2X1 U11880 ( .A(n9638), .B(n2243), .Y(n11690) );
  OR2X1 U11881 ( .A(n9755), .B(n2736), .Y(n12154) );
  OR2X1 U11882 ( .A(n9769), .B(p_1_cast_fu_1031_p1[5]), .Y(n11576) );
  OR2X1 U11883 ( .A(n9501), .B(p_cast_fu_688_p1[5]), .Y(n12209) );
  INVX1 U11884 ( .A(ap_CS_fsm[1]), .Y(n8979) );
  INVX1 U11885 ( .A(ap_CS_fsm[1]), .Y(n8980) );
  OR2X1 U11886 ( .A(n9626), .B(n2251), .Y(n11683) );
  OR2X1 U11887 ( .A(n9741), .B(n2744), .Y(n12147) );
  INVX1 U11888 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/n649 ), 
        .Y(n9469) );
  OR2X1 U11889 ( .A(n9612), .B(n2259), .Y(n11708) );
  OR2X1 U11890 ( .A(n9724), .B(n2752), .Y(n12172) );
  OR2X1 U11891 ( .A(n9598), .B(n2267), .Y(n11701) );
  OR2X1 U11892 ( .A(n9707), .B(n2760), .Y(n12165) );
  OR2X1 U11893 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[0] ), .B(
        n9383), .Y(n8576) );
  OR2X1 U11894 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[0] ), .B(n10205), .Y(n8577) );
  OR2X1 U11895 ( .A(n9707), .B(sum_phi_fu_311_p4[16]), .Y(n11505) );
  OR2X1 U11896 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[2] ), .B(
        n8635), .Y(n8578) );
  OR2X1 U11897 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[2] ), .B(n8634), .Y(n8579) );
  OR2X1 U11898 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[3] ), .B(
        n8578), .Y(n8580) );
  OR2X1 U11899 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[4] ), .B(
        n8580), .Y(n8581) );
  OR2X1 U11900 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[3] ), .B(n8579), .Y(n8582) );
  OR2X1 U11901 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[5] ), .B(
        n8581), .Y(n8583) );
  OR2X1 U11902 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[4] ), .B(n8582), .Y(n8584) );
  OR2X1 U11903 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[6] ), .B(
        n8583), .Y(n8585) );
  OR2X1 U11904 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[5] ), .B(n8584), .Y(n8586) );
  OR2X1 U11905 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[7] ), .B(
        n8585), .Y(n8587) );
  OR2X1 U11906 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[6] ), .B(n8586), .Y(n8588) );
  OR2X1 U11907 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[8] ), .B(
        n8587), .Y(n8589) );
  OR2X1 U11908 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[7] ), .B(n8588), .Y(n8590) );
  OR2X1 U11909 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[9] ), .B(
        n8589), .Y(n8591) );
  OR2X1 U11910 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[8] ), .B(n8590), .Y(n8592) );
  OR2X1 U11911 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[10] ), .B(
        n8591), .Y(n8593) );
  OR2X1 U11912 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[9] ), .B(n8592), .Y(n8594) );
  OR2X1 U11913 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[11] ), .B(
        n8593), .Y(n8595) );
  OR2X1 U11914 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[10] ), .B(n8594), .Y(n8596) );
  OR2X1 U11915 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[12] ), .B(
        n8595), .Y(n8597) );
  OR2X1 U11916 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[11] ), .B(n8596), .Y(n8598) );
  OR2X1 U11917 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[13] ), .B(
        n8597), .Y(n8599) );
  OR2X1 U11918 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[12] ), .B(n8598), .Y(n8600) );
  OR2X1 U11919 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[14] ), .B(
        n8599), .Y(n8601) );
  OR2X1 U11920 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[13] ), .B(n8600), .Y(n8602) );
  OR2X1 U11921 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[15] ), .B(
        n8601), .Y(n8603) );
  OR2X1 U11922 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[14] ), .B(n8602), .Y(n8604) );
  OR2X1 U11923 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[16] ), .B(
        n8603), .Y(n8605) );
  OR2X1 U11924 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[15] ), .B(n8604), .Y(n8606) );
  OR2X1 U11925 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[17] ), .B(
        n8605), .Y(n8607) );
  OR2X1 U11926 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[16] ), .B(n8606), .Y(n8608) );
  OR2X1 U11927 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[18] ), .B(
        n8607), .Y(n8609) );
  OR2X1 U11928 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[17] ), .B(n8608), .Y(n8610) );
  OR2X1 U11929 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[19] ), .B(
        n8609), .Y(n8611) );
  OR2X1 U11930 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[18] ), .B(n8610), .Y(n8612) );
  OR2X1 U11931 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[20] ), .B(
        n8611), .Y(n8613) );
  OR2X1 U11932 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[19] ), .B(n8612), .Y(n8614) );
  OR2X1 U11933 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[21] ), .B(
        n8613), .Y(n8615) );
  OR2X1 U11934 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[20] ), .B(n8614), .Y(n8616) );
  OR2X1 U11935 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[22] ), .B(
        n8615), .Y(n8617) );
  OR2X1 U11936 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[21] ), .B(n8616), .Y(n8618) );
  OR2X1 U11937 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[23] ), .B(
        n8617), .Y(n8619) );
  OR2X1 U11938 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[22] ), .B(n8618), .Y(n8620) );
  OR2X1 U11939 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[24] ), .B(
        n8619), .Y(n8621) );
  OR2X1 U11940 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[23] ), .B(n8620), .Y(n8622) );
  OR2X1 U11941 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[25] ), .B(
        n8621), .Y(n8623) );
  OR2X1 U11942 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[24] ), .B(n8622), .Y(n8624) );
  OR2X1 U11943 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[26] ), .B(
        n8623), .Y(n8625) );
  OR2X1 U11944 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[25] ), .B(n8624), .Y(n8626) );
  OR2X1 U11945 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[27] ), .B(
        n8625), .Y(n8627) );
  OR2X1 U11946 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[26] ), .B(n8626), .Y(n8628) );
  OR2X1 U11947 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[28] ), .B(
        n8627), .Y(n8629) );
  OR2X1 U11948 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[27] ), .B(n8628), .Y(n8630) );
  OR2X1 U11949 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[29] ), .B(
        n8629), .Y(n8631) );
  OR2X1 U11950 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[28] ), .B(n8630), .Y(n8632) );
  OR2X1 U11951 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[29] ), .B(n8632), .Y(n8633) );
  OR2X1 U11952 ( .A(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[1] ), .B(n8577), .Y(n8634) );
  OR2X1 U11953 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[1] ), .B(
        n8576), .Y(n8635) );
  INVX1 U11954 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[25]), .Y(
        n10249) );
  INVX1 U11955 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[21]), .Y(
        n10253) );
  INVX1 U11956 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[25]), .Y(n9941)
         );
  INVX1 U11957 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[21]), .Y(n9945)
         );
  INVX1 U11958 ( .A(p_tmp_i_fu_587_p3[26]), .Y(n9864) );
  INVX1 U11959 ( .A(p_tmp_i_fu_587_p3[22]), .Y(n9868) );
  INVX1 U11960 ( .A(p_tmp_i_fu_587_p3[19]), .Y(n9871) );
  INVX1 U11961 ( .A(p_tmp_i_fu_587_p3[15]), .Y(n9875) );
  AND2X1 U11962 ( .A(n9313), .B(\Decision_AXILiteS_s_axi_U/n248 ), .Y(
        \Decision_AXILiteS_s_axi_U/n155 ) );
  AND2X1 U11963 ( .A(n9312), .B(\Decision_AXILiteS_s_axi_U/n248 ), .Y(
        \Decision_AXILiteS_s_axi_U/n157 ) );
  INVX1 U11964 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[26]), .Y(
        n10248) );
  INVX1 U11965 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[22]), .Y(
        n10252) );
  INVX1 U11966 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[10]), .Y(
        n10264) );
  INVX1 U11967 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[26]), .Y(n9940)
         );
  INVX1 U11968 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[22]), .Y(n9944)
         );
  INVX1 U11969 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[10]), .Y(n9956)
         );
  INVX1 U11970 ( .A(p_tmp_i_fu_587_p3[27]), .Y(n9863) );
  INVX1 U11971 ( .A(p_tmp_i_fu_587_p3[23]), .Y(n9867) );
  INVX1 U11972 ( .A(p_tmp_i_fu_587_p3[16]), .Y(n9874) );
  OR2X1 U11973 ( .A(n9560), .B(n2291), .Y(n11664) );
  OR2X1 U11974 ( .A(n9661), .B(n2784), .Y(n12128) );
  AND2X1 U11975 ( .A(n10901), .B(n10900), .Y(s_axi_AXILiteS_AWREADY) );
  OR2X1 U11976 ( .A(i_8_fu_1148_p2[2]), .B(i_8_fu_1148_p2[1]), .Y(n8638) );
  OR2X1 U11977 ( .A(i_2_fu_823_p2[2]), .B(i_2_fu_823_p2[1]), .Y(n8639) );
  OR2X1 U11978 ( .A(i_11_fu_1179_p2[2]), .B(i_11_fu_1179_p2[1]), .Y(n8640) );
  OR2X1 U11979 ( .A(i_5_fu_854_p2[2]), .B(i_5_fu_854_p2[1]), .Y(n8641) );
  INVX1 U11980 ( .A(n1249), .Y(n10270) );
  AND2X1 U11981 ( .A(tmp_33_i1_fu_1099_p2[2]), .B(tmp_33_i1_fu_1099_p2[1]), 
        .Y(n1250) );
  INVX1 U11982 ( .A(n1811), .Y(n9962) );
  AND2X1 U11983 ( .A(tmp_33_i_fu_786_p2[2]), .B(tmp_33_i_fu_786_p2[1]), .Y(
        n1812) );
  OR2X1 U11984 ( .A(n8922), .B(CircularBuffer_len_read_assign_2_fu_1085_p2[3]), 
        .Y(CircularBuffer_len_read_assign_3_fu_1091_p3[3]) );
  OR2X1 U11985 ( .A(n8920), .B(CircularBuffer_len_read_assign_fu_772_p2[3]), 
        .Y(CircularBuffer_len_read_assign_1_fu_778_p3[3]) );
  INVX1 U11986 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[19]), .Y(
        n10255) );
  INVX1 U11987 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[8]), .Y(n10266) );
  INVX1 U11988 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[19]), .Y(n9947)
         );
  INVX1 U11989 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[8]), .Y(n9958) );
  INVX1 U11990 ( .A(p_tmp_i_fu_587_p3[8]), .Y(n9882) );
  OR2X1 U11991 ( .A(i_8_fu_1148_p2[3]), .B(n8638), .Y(n8642) );
  OR2X1 U11992 ( .A(i_2_fu_823_p2[3]), .B(n8639), .Y(n8643) );
  INVX1 U11993 ( .A(p_tmp_i_fu_587_p3[5]), .Y(n9885) );
  INVX1 U11994 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[20]), .Y(
        n10254) );
  INVX1 U11995 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[9]), .Y(n10265) );
  INVX1 U11996 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[20]), .Y(n9946)
         );
  INVX1 U11997 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[9]), .Y(n9957) );
  INVX1 U11998 ( .A(p_tmp_i_fu_587_p3[10]), .Y(n9880) );
  INVX1 U11999 ( .A(p_tmp_i_fu_587_p3[9]), .Y(n9881) );
  INVX1 U12000 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[18]), .Y(n9948)
         );
  INVX1 U12001 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[7]), .Y(n9959) );
  INVX1 U12002 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[18]), .Y(
        n10256) );
  INVX1 U12003 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[7]), .Y(n10267) );
  INVX1 U12004 ( .A(p_tmp_i_fu_587_p3[7]), .Y(n9883) );
  INVX1 U12005 ( .A(\Decision_AXILiteS_s_axi_U/n630 ), .Y(n8918) );
  AND2X1 U12006 ( .A(n11495), .B(n9661), .Y(n11496) );
  AND2X1 U12007 ( .A(n11790), .B(n9598), .Y(n11791) );
  AND2X1 U12008 ( .A(n11797), .B(n9612), .Y(n11798) );
  AND2X1 U12009 ( .A(n11532), .B(n9707), .Y(n11533) );
  AND2X1 U12010 ( .A(n10899), .B(n10898), .Y(\Decision_AXILiteS_s_axi_U/n575 )
         );
  INVX1 U12011 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[17]), .Y(n9949)
         );
  INVX1 U12012 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[6]), .Y(n9960) );
  INVX1 U12013 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[17]), .Y(
        n10257) );
  INVX1 U12014 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[6]), .Y(n10268) );
  INVX1 U12015 ( .A(p_tmp_i_fu_587_p3[6]), .Y(n9884) );
  AND2X1 U12016 ( .A(n11162), .B(n10719), .Y(n11163) );
  INVX1 U12017 ( .A(ap_CS_fsm[4]), .Y(n9011) );
  AND2X1 U12018 ( .A(n11664), .B(n9558), .Y(n11665) );
  AND2X1 U12019 ( .A(n12128), .B(n9659), .Y(n12129) );
  INVX1 U12020 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[5]), .Y(n9961) );
  INVX1 U12021 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[5]), .Y(n10269) );
  INVX1 U12022 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[14]), .Y(n9952)
         );
  INVX1 U12023 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[16]), .Y(n9950)
         );
  INVX1 U12024 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[12]), .Y(n9954)
         );
  INVX1 U12025 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[30]), .Y(n9936)
         );
  INVX1 U12026 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[28]), .Y(n9938)
         );
  INVX1 U12027 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[24]), .Y(n9942)
         );
  INVX1 U12028 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[30]), .Y(
        n10244) );
  INVX1 U12029 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[28]), .Y(
        n10246) );
  INVX1 U12030 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[24]), .Y(
        n10250) );
  INVX1 U12031 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[16]), .Y(
        n10258) );
  INVX1 U12032 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[14]), .Y(
        n10260) );
  INVX1 U12033 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[12]), .Y(
        n10262) );
  INVX1 U12034 ( .A(p_tmp_i_fu_587_p3[12]), .Y(n9878) );
  INVX1 U12035 ( .A(p_tmp_i_fu_587_p3[14]), .Y(n9876) );
  INVX1 U12036 ( .A(p_tmp_i_fu_587_p3[18]), .Y(n9872) );
  INVX1 U12037 ( .A(p_tmp_i_fu_587_p3[21]), .Y(n9869) );
  INVX1 U12038 ( .A(p_tmp_i_fu_587_p3[25]), .Y(n9865) );
  INVX1 U12039 ( .A(p_tmp_i_fu_587_p3[29]), .Y(n9861) );
  AND2X1 U12040 ( .A(n11701), .B(n9596), .Y(n11702) );
  AND2X1 U12041 ( .A(n12165), .B(n9705), .Y(n12166) );
  AND2X1 U12042 ( .A(n12076), .B(n9705), .Y(n12077) );
  AND2X1 U12043 ( .A(n12083), .B(n9721), .Y(n12084) );
  AND2X1 U12044 ( .A(n11987), .B(n9596), .Y(n11988) );
  AND2X1 U12045 ( .A(n11994), .B(n9610), .Y(n11995) );
  INVX1 U12046 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[13]), .Y(n9953)
         );
  INVX1 U12047 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[15]), .Y(n9951)
         );
  INVX1 U12048 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[11]), .Y(n9955)
         );
  INVX1 U12049 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[29]), .Y(n9937)
         );
  INVX1 U12050 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[27]), .Y(n9939)
         );
  INVX1 U12051 ( .A(CircularBuffer_head_i_read_ass_fu_797_p3[23]), .Y(n9943)
         );
  INVX1 U12052 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[29]), .Y(
        n10245) );
  INVX1 U12053 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[27]), .Y(
        n10247) );
  INVX1 U12054 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[23]), .Y(
        n10251) );
  INVX1 U12055 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[15]), .Y(
        n10259) );
  INVX1 U12056 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[13]), .Y(
        n10261) );
  INVX1 U12057 ( .A(CircularBuffer_head_i_read_ass_1_fu_1110_p3[11]), .Y(
        n10263) );
  INVX1 U12058 ( .A(p_tmp_i_fu_587_p3[11]), .Y(n9879) );
  INVX1 U12059 ( .A(p_tmp_i_fu_587_p3[13]), .Y(n9877) );
  INVX1 U12060 ( .A(p_tmp_i_fu_587_p3[17]), .Y(n9873) );
  INVX1 U12061 ( .A(p_tmp_i_fu_587_p3[20]), .Y(n9870) );
  INVX1 U12062 ( .A(p_tmp_i_fu_587_p3[24]), .Y(n9866) );
  INVX1 U12063 ( .A(p_tmp_i_fu_587_p3[28]), .Y(n9862) );
  INVX1 U12064 ( .A(p_tmp_i_fu_587_p3[30]), .Y(n9860) );
  AND2X1 U12065 ( .A(n11155), .B(n10711), .Y(n11156) );
  AND2X1 U12066 ( .A(n11879), .B(n10409), .Y(n11880) );
  AND2X1 U12067 ( .A(n11886), .B(n10420), .Y(n11887) );
  INVX1 U12068 ( .A(ap_rst_n), .Y(n9042) );
  OR2X1 U12069 ( .A(n9596), .B(n2269), .Y(n11674) );
  OR2X1 U12070 ( .A(n9705), .B(n2762), .Y(n12138) );
  INVX1 U12071 ( .A(\reset_V_V[0] ), .Y(n8897) );
  INVX1 U12072 ( .A(\reset_A_V[0] ), .Y(n8898) );
  INVX1 U12073 ( .A(n8872), .Y(n10058) );
  INVX1 U12074 ( .A(n8871), .Y(n10059) );
  INVX1 U12075 ( .A(n8875), .Y(n9930) );
  INVX1 U12076 ( .A(n8874), .Y(n9931) );
  INVX1 U12077 ( .A(n8870), .Y(n10060) );
  INVX1 U12078 ( .A(n8873), .Y(n9932) );
  AND2X1 U12079 ( .A(n10896), .B(\Decision_AXILiteS_s_axi_U/waddr[3] ), .Y(
        \Decision_AXILiteS_s_axi_U/n611 ) );
  INVX1 U12080 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[24]), .Y(n9336) );
  INVX1 U12081 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[24]), .Y(n10180) );
  INVX1 U12082 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[6]), .Y(n9373)
         );
  INVX1 U12083 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[2]), .Y(n9379)
         );
  INVX1 U12084 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[10]), .Y(n9365) );
  INVX1 U12085 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[14]), .Y(n9358) );
  INVX1 U12086 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[18]), .Y(n9349) );
  INVX1 U12087 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[22]), .Y(n9342) );
  INVX1 U12088 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[10]), .Y(n10194) );
  INVX1 U12089 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[14]), .Y(n10190) );
  INVX1 U12090 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[18]), .Y(n10186) );
  INVX1 U12091 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[22]), .Y(n10182) );
  INVX1 U12092 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[26]), .Y(n10178) );
  INVX1 U12093 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[26]), .Y(n9334) );
  INVX1 U12094 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[6]), .Y(n10198)
         );
  INVX1 U12095 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[2]), .Y(n10202)
         );
  INVX1 U12096 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[4]), .Y(n9375)
         );
  INVX1 U12097 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[4]), .Y(n10200)
         );
  INVX1 U12098 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[1]), .Y(n9381)
         );
  INVX1 U12099 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[1]), .Y(n10203)
         );
  INVX1 U12100 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[12]), .Y(n9360) );
  INVX1 U12101 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[12]), .Y(n10192) );
  INVX1 U12102 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[28]), .Y(n10176) );
  INVX1 U12103 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[28]), .Y(n9329) );
  INVX1 U12104 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[16]), .Y(n9351) );
  INVX1 U12105 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[20]), .Y(n9344) );
  INVX1 U12106 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[16]), .Y(n10188) );
  INVX1 U12107 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[20]), .Y(n10184) );
  INVX1 U12108 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[5]), .Y(n9374)
         );
  INVX1 U12109 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[21]), .Y(n10183) );
  INVX1 U12110 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[17]), .Y(n9350) );
  INVX1 U12111 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[21]), .Y(n9343) );
  INVX1 U12112 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[17]), .Y(n10187) );
  INVX1 U12113 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[5]), .Y(n10199)
         );
  INVX1 U12114 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[31]), .Y(n10173) );
  INVX1 U12115 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[31]), .Y(n9326) );
  INVX1 U12116 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[30]), .Y(n10174) );
  INVX1 U12117 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[30]), .Y(n9327) );
  INVX1 U12118 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[9]), .Y(n9367)
         );
  INVX1 U12119 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[9]), .Y(n10195)
         );
  INVX1 U12120 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[13]), .Y(n9359) );
  INVX1 U12121 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[13]), .Y(n10191) );
  INVX1 U12122 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[29]), .Y(n10175) );
  INVX1 U12123 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[25]), .Y(n10179) );
  INVX1 U12124 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[29]), .Y(n9328) );
  INVX1 U12125 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[25]), .Y(n9335) );
  INVX1 U12126 ( .A(sum_1_phi_fu_379_p4[31]), .Y(n9325) );
  INVX1 U12127 ( .A(sum_phi_fu_311_p4[31]), .Y(n10070) );
  INVX1 U12128 ( .A(n7853), .Y(n10301) );
  INVX1 U12129 ( .A(n7634), .Y(n10019) );
  INVX1 U12130 ( .A(n7636), .Y(n10328) );
  INVX1 U12131 ( .A(n7851), .Y(n9987) );
  INVX1 U12132 ( .A(n11267), .Y(n10299) );
  INVX1 U12133 ( .A(n11371), .Y(n10017) );
  INVX1 U12134 ( .A(n11423), .Y(n10326) );
  INVX1 U12135 ( .A(n11319), .Y(n9985) );
  INVX1 U12136 ( .A(n11271), .Y(n10297) );
  INVX1 U12137 ( .A(n11375), .Y(n10015) );
  INVX1 U12138 ( .A(n11427), .Y(n10324) );
  INVX1 U12139 ( .A(n11323), .Y(n9983) );
  INVX1 U12140 ( .A(n11275), .Y(n10295) );
  INVX1 U12141 ( .A(n11379), .Y(n10013) );
  INVX1 U12142 ( .A(n11431), .Y(n10322) );
  INVX1 U12143 ( .A(n11327), .Y(n9981) );
  INVX1 U12144 ( .A(n11279), .Y(n10293) );
  INVX1 U12145 ( .A(n11383), .Y(n10011) );
  INVX1 U12146 ( .A(n11435), .Y(n10320) );
  INVX1 U12147 ( .A(n11331), .Y(n9979) );
  INVX1 U12148 ( .A(n11283), .Y(n10291) );
  INVX1 U12149 ( .A(n11387), .Y(n10009) );
  INVX1 U12150 ( .A(n11439), .Y(n10318) );
  INVX1 U12151 ( .A(n11335), .Y(n9977) );
  INVX1 U12152 ( .A(n11287), .Y(n10289) );
  INVX1 U12153 ( .A(n11391), .Y(n10007) );
  INVX1 U12154 ( .A(n11443), .Y(n10316) );
  INVX1 U12155 ( .A(n11339), .Y(n9975) );
  INVX1 U12156 ( .A(n11291), .Y(n10287) );
  INVX1 U12157 ( .A(n11395), .Y(n10005) );
  INVX1 U12158 ( .A(n11447), .Y(n10314) );
  INVX1 U12159 ( .A(n11343), .Y(n9973) );
  INVX1 U12160 ( .A(n11295), .Y(n10285) );
  INVX1 U12161 ( .A(n11399), .Y(n10003) );
  INVX1 U12162 ( .A(n11451), .Y(n10312) );
  INVX1 U12163 ( .A(n11347), .Y(n9971) );
  INVX1 U12164 ( .A(n11299), .Y(n10283) );
  INVX1 U12165 ( .A(n11403), .Y(n10001) );
  INVX1 U12166 ( .A(n8093), .Y(n10310) );
  INVX1 U12167 ( .A(n8091), .Y(n9969) );
  INVX1 U12168 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[0]), .Y(n9382)
         );
  INVX1 U12169 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[0]), .Y(n10204)
         );
  INVX1 U12170 ( .A(n8644), .Y(recentVBools_data_address0[1]) );
  OR2X1 U12171 ( .A(p_tmp_i_reg_1556[29]), .B(p_tmp_i_reg_1556[28]), .Y(n11236) );
  INVX1 U12172 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[7]), .Y(n9372)
         );
  INVX1 U12173 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[3]), .Y(n9378)
         );
  INVX1 U12174 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[8]), .Y(n9369)
         );
  INVX1 U12175 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[11]), .Y(n9364) );
  INVX1 U12176 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[15]), .Y(n9357) );
  INVX1 U12177 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[11]), .Y(n10193) );
  INVX1 U12178 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[15]), .Y(n10189) );
  INVX1 U12179 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[23]), .Y(n10181) );
  INVX1 U12180 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[19]), .Y(n9348) );
  INVX1 U12181 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[7]), .Y(n10197)
         );
  INVX1 U12182 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[27]), .Y(n10177) );
  INVX1 U12183 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[19]), .Y(n10185) );
  INVX1 U12184 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[27]), .Y(n9333) );
  INVX1 U12185 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[3]), .Y(n10201)
         );
  INVX1 U12186 ( .A(CircularBuffer_sum_write_assig_1_fu_917_p2[8]), .Y(n10196)
         );
  INVX1 U12187 ( .A(CircularBuffer_sum_write_assig_3_fu_1242_p2[23]), .Y(n9341) );
  OR2X1 U12188 ( .A(n9753), .B(tmp_7_reg_1544[28]), .Y(n12053) );
  OR2X1 U12189 ( .A(n9636), .B(tmp_6_reg_1538[28]), .Y(n11964) );
  OR2X1 U12190 ( .A(n10441), .B(VbeatDelay_new_1_reg_326[28]), .Y(n11856) );
  OR2X1 U12191 ( .A(n10735), .B(VbeatDelay_new_1_reg_326[28]), .Y(n11132) );
  BUFX2 U12192 ( .A(recentdatapoints_data_address0[0]), .Y(n8888) );
  OR2X1 U12193 ( .A(n9690), .B(tmp_7_reg_1544[12]), .Y(n12008) );
  OR2X1 U12194 ( .A(n9584), .B(tmp_6_reg_1538[12]), .Y(n11919) );
  OR2X1 U12195 ( .A(n10399), .B(VbeatDelay_new_1_reg_326[12]), .Y(n11811) );
  OR2X1 U12196 ( .A(n10703), .B(VbeatDelay_new_1_reg_326[12]), .Y(n11087) );
  INVX1 U12197 ( .A(n8645), .Y(recentABools_data_address0[1]) );
  OR2X1 U12198 ( .A(VbeatFallDelay_new_1_reg_342[26]), .B(
        VbeatFallDelay_new_1_reg_342[25]), .Y(n11899) );
  INVX1 U12199 ( .A(a_thresh[20]), .Y(n9780) );
  INVX1 U12200 ( .A(a_thresh[23]), .Y(n9783) );
  INVX1 U12201 ( .A(a_thresh[18]), .Y(n9778) );
  INVX1 U12202 ( .A(v_thresh[20]), .Y(n9521) );
  INVX1 U12203 ( .A(v_thresh[23]), .Y(n9524) );
  INVX1 U12204 ( .A(v_thresh[18]), .Y(n9519) );
  OR2X1 U12205 ( .A(AbeatDelay_new_reg_394[30]), .B(AbeatDelay_new_reg_394[29]), .Y(n11050) );
  OR2X1 U12206 ( .A(AbeatDelay_new_reg_394[30]), .B(AbeatDelay_new_reg_394[29]), .Y(n11070) );
  OR2X1 U12207 ( .A(AbeatDelay_new_reg_394[26]), .B(AbeatDelay_new_reg_394[25]), .Y(n11049) );
  OR2X1 U12208 ( .A(AbeatDelay_new_reg_394[26]), .B(AbeatDelay_new_reg_394[25]), .Y(n11069) );
  INVX1 U12209 ( .A(ap_start), .Y(n10889) );
  INVX1 U12210 ( .A(n11085), .Y(n10674) );
  AND2X1 U12211 ( .A(n12039), .B(n9659), .Y(n12040) );
  AND2X1 U12212 ( .A(n11950), .B(n9558), .Y(n11951) );
  INVX1 U12213 ( .A(sum_1_phi_fu_379_p4[1]), .Y(n9380) );
  INVX1 U12214 ( .A(n11154), .Y(n10498) );
  INVX1 U12215 ( .A(n11700), .Y(n9601) );
  INVX1 U12216 ( .A(n12164), .Y(n9712) );
  INVX1 U12217 ( .A(n12075), .Y(n9710) );
  INVX1 U12218 ( .A(n11986), .Y(n9603) );
  INVX1 U12219 ( .A(n11878), .Y(n10414) );
  INVX1 U12220 ( .A(n11789), .Y(n9346) );
  INVX1 U12221 ( .A(n11531), .Y(n9716) );
  AND2X1 U12222 ( .A(n11842), .B(n10377), .Y(n11843) );
  AND2X1 U12223 ( .A(n11118), .B(n10686), .Y(n11119) );
  INVX1 U12224 ( .A(a_thresh[17]), .Y(n9777) );
  INVX1 U12225 ( .A(a_thresh[16]), .Y(n9776) );
  INVX1 U12226 ( .A(v_thresh[17]), .Y(n9518) );
  INVX1 U12227 ( .A(v_thresh[16]), .Y(n9517) );
  INVX1 U12228 ( .A(n2195), .Y(n10278) );
  INVX1 U12229 ( .A(n2201), .Y(n9996) );
  OR2X1 U12230 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[0]), .B(n10634), 
        .Y(n8646) );
  OR2X1 U12231 ( .A(CircularBuffer_head_i_read_ass_reg_1624[0]), .B(n10139), 
        .Y(n8647) );
  OR2X1 U12232 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[0]), .B(n10541), 
        .Y(n8648) );
  OR2X1 U12233 ( .A(CircularBuffer_head_i_read_ass_reg_1624[0]), .B(n10076), 
        .Y(n8649) );
  INVX1 U12234 ( .A(n11161), .Y(n10509) );
  INVX1 U12235 ( .A(n11494), .Y(n9667) );
  INVX1 U12236 ( .A(n11663), .Y(n9562) );
  INVX1 U12237 ( .A(n12127), .Y(n9664) );
  INVX1 U12238 ( .A(n12082), .Y(n9727) );
  INVX1 U12239 ( .A(n11993), .Y(n9617) );
  INVX1 U12240 ( .A(n11885), .Y(n10425) );
  INVX1 U12241 ( .A(n11796), .Y(n9339) );
  BUFX2 U12242 ( .A(recentdatapoints_data_address0[1]), .Y(n8889) );
  INVX1 U12243 ( .A(CircularBuffer_len_read_assign_3_reg_1711[1]), .Y(n10574)
         );
  INVX1 U12244 ( .A(CircularBuffer_len_read_assign_1_reg_1616[1]), .Y(n10079)
         );
  INVX1 U12245 ( .A(n11067), .Y(n10673) );
  INVX1 U12246 ( .A(a_thresh[1]), .Y(n9766) );
  INVX1 U12247 ( .A(v_thresh[1]), .Y(n9497) );
  INVX1 U12248 ( .A(a_thresh[25]), .Y(n9785) );
  INVX1 U12249 ( .A(a_thresh[24]), .Y(n9784) );
  INVX1 U12250 ( .A(v_thresh[25]), .Y(n9527) );
  INVX1 U12251 ( .A(v_thresh[24]), .Y(n9526) );
  INVX1 U12252 ( .A(a_thresh[26]), .Y(n9786) );
  INVX1 U12253 ( .A(v_thresh[26]), .Y(n9528) );
  INVX1 U12254 ( .A(\not_tmp_i_i2_reg_1745[0] ), .Y(n10668) );
  INVX1 U12255 ( .A(\not_tmp_i_i4_reg_1650[0] ), .Y(n10171) );
  INVX1 U12256 ( .A(n11077), .Y(n10676) );
  INVX1 U12257 ( .A(n11411), .Y(n10331) );
  INVX1 U12258 ( .A(n11307), .Y(n9990) );
  INVX1 U12259 ( .A(n8098), .Y(n10281) );
  INVX1 U12260 ( .A(n7850), .Y(n9999) );
  INVX1 U12261 ( .A(n8368), .Y(n10308) );
  INVX1 U12262 ( .A(n8365), .Y(n9967) );
  INVX1 U12263 ( .A(n11255), .Y(n10304) );
  INVX1 U12264 ( .A(n11359), .Y(n10022) );
  AND2X1 U12265 ( .A(ap_rst_n), .B(n5294), .Y(n8650) );
  INVX1 U12266 ( .A(n8650), .Y(\Decision_AXILiteS_s_axi_U/n533 ) );
  AND2X1 U12267 ( .A(ap_rst_n), .B(n5293), .Y(n8651) );
  INVX1 U12268 ( .A(n8651), .Y(\Decision_AXILiteS_s_axi_U/n429 ) );
  INVX1 U12269 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[15] ), .Y(n10883)
         );
  INVX1 U12270 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[14] ), .Y(n10882)
         );
  INVX1 U12271 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[13] ), .Y(n10881)
         );
  INVX1 U12272 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[12] ), .Y(n10880)
         );
  INVX1 U12273 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[11] ), .Y(n10879)
         );
  INVX1 U12274 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[10] ), .Y(n10878)
         );
  INVX1 U12275 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[9] ), .Y(n10877)
         );
  INVX1 U12276 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[8] ), .Y(n10876)
         );
  INVX1 U12277 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[7] ), .Y(n10875)
         );
  INVX1 U12278 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[6] ), .Y(n10874)
         );
  INVX1 U12279 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[5] ), .Y(n10873)
         );
  INVX1 U12280 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[4] ), .Y(n10872)
         );
  INVX1 U12281 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[3] ), .Y(n10871)
         );
  INVX1 U12282 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[2] ), .Y(n10870)
         );
  INVX1 U12283 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[1] ), .Y(n10869)
         );
  INVX1 U12284 ( .A(\Decision_AXILiteS_s_axi_U/int_ap_return[0] ), .Y(n10868)
         );
  INVX1 U12285 ( .A(CircularBuffer_len_read_assign_3_reg_1711[10]), .Y(n10583)
         );
  INVX1 U12286 ( .A(CircularBuffer_len_read_assign_3_reg_1711[9]), .Y(n10582)
         );
  INVX1 U12287 ( .A(CircularBuffer_len_read_assign_3_reg_1711[8]), .Y(n10581)
         );
  INVX1 U12288 ( .A(\tmp_13_reg_1725[0] ), .Y(n10542) );
  INVX1 U12289 ( .A(recentABools_head_i[1]), .Y(n10363) );
  INVX1 U12290 ( .A(CircularBuffer_len_read_assign_3_reg_1711[23]), .Y(n10596)
         );
  INVX1 U12291 ( .A(CircularBuffer_len_read_assign_3_reg_1711[22]), .Y(n10595)
         );
  INVX1 U12292 ( .A(CircularBuffer_len_read_assign_3_reg_1711[14]), .Y(n10587)
         );
  INVX1 U12293 ( .A(CircularBuffer_len_read_assign_3_reg_1711[13]), .Y(n10586)
         );
  INVX1 U12294 ( .A(recentABools_head_i[2]), .Y(n10361) );
  INVX1 U12295 ( .A(recentABools_head_i[3]), .Y(n10359) );
  INVX1 U12296 ( .A(recentABools_head_i[4]), .Y(n10357) );
  INVX1 U12297 ( .A(CircularBuffer_len_read_assign_3_reg_1711[29]), .Y(n10602)
         );
  INVX1 U12298 ( .A(CircularBuffer_len_read_assign_3_reg_1711[28]), .Y(n10601)
         );
  INVX1 U12299 ( .A(CircularBuffer_len_read_assign_3_reg_1711[25]), .Y(n10598)
         );
  INVX1 U12300 ( .A(CircularBuffer_len_read_assign_3_reg_1711[24]), .Y(n10597)
         );
  INVX1 U12301 ( .A(AbeatDelay_new_reg_394[27]), .Y(n10733) );
  INVX1 U12302 ( .A(AbeatDelay_new_reg_394[23]), .Y(n10725) );
  INVX1 U12303 ( .A(AbeatDelay_new_reg_394[19]), .Y(n10717) );
  INVX1 U12304 ( .A(AbeatDelay_new_reg_394[15]), .Y(n10709) );
  INVX1 U12305 ( .A(AbeatDelay_new_reg_394[11]), .Y(n10701) );
  INVX1 U12306 ( .A(AbeatDelay_new_reg_394[3]), .Y(n10683) );
  INVX1 U12307 ( .A(\Decision_AXILiteS_s_axi_U/int_ier[1] ), .Y(n10887) );
  INVX1 U12308 ( .A(recentABools_len[26]), .Y(n10630) );
  INVX1 U12309 ( .A(recentABools_len[25]), .Y(n10629) );
  INVX1 U12310 ( .A(recentABools_len[22]), .Y(n10626) );
  INVX1 U12311 ( .A(recentABools_len[21]), .Y(n10625) );
  INVX1 U12312 ( .A(recentABools_len[20]), .Y(n10624) );
  INVX1 U12313 ( .A(recentABools_len[19]), .Y(n10623) );
  INVX1 U12314 ( .A(recentABools_len[10]), .Y(n10614) );
  INVX1 U12315 ( .A(recentABools_len[9]), .Y(n10613) );
  INVX1 U12316 ( .A(recentABools_len[8]), .Y(n10612) );
  INVX1 U12317 ( .A(recentABools_len[2]), .Y(n10606) );
  INVX1 U12318 ( .A(recentABools_len[1]), .Y(n10605) );
  INVX1 U12319 ( .A(recentABools_data_addr_reg_1689[1]), .Y(n10364) );
  INVX1 U12320 ( .A(recentABools_data_addr_reg_1689[2]), .Y(n10362) );
  INVX1 U12321 ( .A(recentABools_data_addr_reg_1689[3]), .Y(n10360) );
  INVX1 U12322 ( .A(recentABools_data_addr_reg_1689[4]), .Y(n10358) );
  INVX1 U12323 ( .A(recentABools_data_addr_reg_1689[0]), .Y(n10272) );
  INVX1 U12324 ( .A(\last_sample_is_V_V_loc_2_reg_358[0] ), .Y(n10239) );
  INVX1 U12325 ( .A(recentVBools_len[10]), .Y(n10119) );
  INVX1 U12326 ( .A(recentVBools_len[9]), .Y(n10118) );
  INVX1 U12327 ( .A(recentVBools_len[8]), .Y(n10117) );
  INVX1 U12328 ( .A(recentVBools_len[2]), .Y(n10111) );
  INVX1 U12329 ( .A(recentVBools_len[1]), .Y(n10110) );
  INVX1 U12330 ( .A(\Decision_AXILiteS_s_axi_U/int_auto_restart ), .Y(n10890)
         );
  INVX1 U12331 ( .A(recentVBools_len[26]), .Y(n10135) );
  INVX1 U12332 ( .A(recentVBools_len[25]), .Y(n10134) );
  INVX1 U12333 ( .A(recentVBools_len[22]), .Y(n10131) );
  INVX1 U12334 ( .A(recentVBools_len[21]), .Y(n10130) );
  INVX1 U12335 ( .A(recentVBools_len[20]), .Y(n10129) );
  INVX1 U12336 ( .A(recentVBools_len[19]), .Y(n10128) );
  INVX1 U12337 ( .A(VbeatDelay_new_1_reg_326[28]), .Y(n10525) );
  INVX1 U12338 ( .A(VbeatDelay_new_1_reg_326[24]), .Y(n10515) );
  INVX1 U12339 ( .A(VbeatDelay_new_1_reg_326[20]), .Y(n10504) );
  INVX1 U12340 ( .A(VbeatDelay_new_1_reg_326[17]), .Y(n10495) );
  INVX1 U12341 ( .A(VbeatDelay_new_1_reg_326[16]), .Y(n10493) );
  INVX1 U12342 ( .A(VbeatDelay_new_1_reg_326[10]), .Y(n10478) );
  INVX1 U12343 ( .A(VbeatDelay_new_1_reg_326[4]), .Y(n10461) );
  INVX1 U12344 ( .A(VbeatFallDelay_new_1_reg_342[27]), .Y(n10439) );
  INVX1 U12345 ( .A(VbeatFallDelay_new_1_reg_342[23]), .Y(n10428) );
  INVX1 U12346 ( .A(VbeatFallDelay_new_1_reg_342[19]), .Y(n10417) );
  INVX1 U12347 ( .A(VbeatFallDelay_new_1_reg_342[15]), .Y(n10407) );
  INVX1 U12348 ( .A(VbeatFallDelay_new_1_reg_342[11]), .Y(n10396) );
  INVX1 U12349 ( .A(VbeatFallDelay_new_1_reg_342[8]), .Y(n10388) );
  INVX1 U12350 ( .A(VbeatFallDelay_new_1_reg_342[7]), .Y(n10384) );
  INVX1 U12351 ( .A(VbeatFallDelay_new_1_reg_342[3]), .Y(n10375) );
  INVX1 U12352 ( .A(VbeatFallDelay_new_1_reg_342[0]), .Y(n10368) );
  INVX1 U12353 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][15] ), .Y(n11045) );
  INVX1 U12354 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][14] ), .Y(n11044) );
  INVX1 U12355 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][13] ), .Y(n11043) );
  INVX1 U12356 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][12] ), .Y(n11042) );
  INVX1 U12357 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][7] ), .Y(n11037) );
  INVX1 U12358 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][6] ), .Y(n11036) );
  INVX1 U12359 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][5] ), .Y(n11035) );
  INVX1 U12360 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][4] ), .Y(n11034) );
  INVX1 U12361 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][3] ), .Y(n11033) );
  INVX1 U12362 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][2] ), .Y(n11032) );
  INVX1 U12363 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][1] ), .Y(n11031) );
  INVX1 U12364 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][0] ), .Y(n11030) );
  INVX1 U12365 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][11] ), .Y(n11041) );
  INVX1 U12366 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][10] ), .Y(n11040) );
  INVX1 U12367 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][9] ), .Y(n11039) );
  INVX1 U12368 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[19][8] ), .Y(n11038) );
  INVX1 U12369 ( .A(\last_sample_is_A_V[0] ), .Y(n10810) );
  INVX1 U12370 ( .A(\tmp_25_reg_1777[0] ), .Y(n10809) );
  INVX1 U12371 ( .A(\tmp_22_reg_1772[0] ), .Y(n10775) );
  INVX1 U12372 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][15] ), .Y(n10917) );
  INVX1 U12373 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][14] ), .Y(n10916) );
  INVX1 U12374 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][13] ), .Y(n10915) );
  INVX1 U12375 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][12] ), .Y(n10914) );
  INVX1 U12376 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][7] ), .Y(n10909) );
  INVX1 U12377 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][6] ), .Y(n10908) );
  INVX1 U12378 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][5] ), .Y(n10907) );
  INVX1 U12379 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][4] ), .Y(n10906) );
  INVX1 U12380 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][3] ), .Y(n10905) );
  INVX1 U12381 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][2] ), .Y(n10904) );
  INVX1 U12382 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][1] ), .Y(n10903) );
  INVX1 U12383 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][0] ), .Y(n10902) );
  INVX1 U12384 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][11] ), .Y(n10913) );
  INVX1 U12385 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][10] ), .Y(n10912) );
  INVX1 U12386 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][9] ), .Y(n10911) );
  INVX1 U12387 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[0][8] ), .Y(n10910) );
  INVX1 U12388 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][15] ), .Y(n10965) );
  INVX1 U12389 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][14] ), .Y(n10964) );
  INVX1 U12390 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][13] ), .Y(n10963) );
  INVX1 U12391 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][12] ), .Y(n10962) );
  INVX1 U12392 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][7] ), .Y(n10957) );
  INVX1 U12393 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][6] ), .Y(n10956) );
  INVX1 U12394 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][5] ), .Y(n10955) );
  INVX1 U12395 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][4] ), .Y(n10954) );
  INVX1 U12396 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][3] ), .Y(n10953) );
  INVX1 U12397 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][2] ), .Y(n10952) );
  INVX1 U12398 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][1] ), .Y(n10951) );
  INVX1 U12399 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][0] ), .Y(n10950) );
  INVX1 U12400 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][15] ), .Y(n10933) );
  INVX1 U12401 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][14] ), .Y(n10932) );
  INVX1 U12402 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][13] ), .Y(n10931) );
  INVX1 U12403 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][12] ), .Y(n10930) );
  INVX1 U12404 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][7] ), .Y(n10925) );
  INVX1 U12405 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][6] ), .Y(n10924) );
  INVX1 U12406 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][5] ), .Y(n10923) );
  INVX1 U12407 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][4] ), .Y(n10922) );
  INVX1 U12408 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][3] ), .Y(n10921) );
  INVX1 U12409 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][2] ), .Y(n10920) );
  INVX1 U12410 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][1] ), .Y(n10919) );
  INVX1 U12411 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][0] ), .Y(n10918) );
  INVX1 U12412 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][11] ), .Y(n10961) );
  INVX1 U12413 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][10] ), .Y(n10960) );
  INVX1 U12414 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][9] ), .Y(n10959) );
  INVX1 U12415 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[3][8] ), .Y(n10958) );
  INVX1 U12416 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][15] ), .Y(n10949) );
  INVX1 U12417 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][14] ), .Y(n10948) );
  INVX1 U12418 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][13] ), .Y(n10947) );
  INVX1 U12419 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][12] ), .Y(n10946) );
  INVX1 U12420 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][7] ), .Y(n10941) );
  INVX1 U12421 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][6] ), .Y(n10940) );
  INVX1 U12422 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][5] ), .Y(n10939) );
  INVX1 U12423 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][4] ), .Y(n10938) );
  INVX1 U12424 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][3] ), .Y(n10937) );
  INVX1 U12425 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][2] ), .Y(n10936) );
  INVX1 U12426 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][1] ), .Y(n10935) );
  INVX1 U12427 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][0] ), .Y(n10934) );
  INVX1 U12428 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][11] ), .Y(n10929) );
  INVX1 U12429 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][10] ), .Y(n10928) );
  INVX1 U12430 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][9] ), .Y(n10927) );
  INVX1 U12431 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[1][8] ), .Y(n10926) );
  INVX1 U12432 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][11] ), .Y(n10945) );
  INVX1 U12433 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][10] ), .Y(n10944) );
  INVX1 U12434 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][9] ), .Y(n10943) );
  INVX1 U12435 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[2][8] ), .Y(n10942) );
  AND2X1 U12436 ( .A(VstimDelay[31]), .B(n8897), .Y(\dp_cluster_0/N985 ) );
  AND2X1 U12437 ( .A(AstimDelay[31]), .B(n8898), .Y(\dp_cluster_1/N953 ) );
  INVX1 U12438 ( .A(recentdatapoints_data_addr_reg_1533[2]), .Y(n9895) );
  INVX1 U12439 ( .A(recentdatapoints_data_addr_reg_1533[3]), .Y(n9891) );
  INVX1 U12440 ( .A(VCaptureThresh[24]), .Y(n9735) );
  INVX1 U12441 ( .A(VCaptureThresh[23]), .Y(n9731) );
  INVX1 U12442 ( .A(VCaptureThresh[22]), .Y(n9725) );
  INVX1 U12443 ( .A(VCaptureThresh[21]), .Y(n9722) );
  INVX1 U12444 ( .A(VCaptureThresh[20]), .Y(n9718) );
  INVX1 U12445 ( .A(VCaptureThresh[19]), .Y(n9714) );
  INVX1 U12446 ( .A(VCaptureThresh[18]), .Y(n9708) );
  INVX1 U12447 ( .A(VCaptureThresh[17]), .Y(n9706) );
  INVX1 U12448 ( .A(VCaptureThresh[16]), .Y(n9704) );
  INVX1 U12449 ( .A(VCaptureThresh[15]), .Y(n9700) );
  INVX1 U12450 ( .A(VCaptureThresh[14]), .Y(n9694) );
  INVX1 U12451 ( .A(VCaptureThresh[13]), .Y(n9691) );
  INVX1 U12452 ( .A(VCaptureThresh[12]), .Y(n9688) );
  INVX1 U12453 ( .A(VCaptureThresh[11]), .Y(n9684) );
  INVX1 U12454 ( .A(VCaptureThresh[10]), .Y(n9678) );
  INVX1 U12455 ( .A(VCaptureThresh[9]), .Y(n9674) );
  INVX1 U12456 ( .A(VCaptureThresh[8]), .Y(n9669) );
  INVX1 U12457 ( .A(VCaptureThresh[7]), .Y(n9666) );
  INVX1 U12458 ( .A(VCaptureThresh[6]), .Y(n9662) );
  INVX1 U12459 ( .A(VCaptureThresh[5]), .Y(n9660) );
  INVX1 U12460 ( .A(VCaptureThresh[4]), .Y(n9658) );
  INVX1 U12461 ( .A(VCaptureThresh[3]), .Y(n9655) );
  INVX1 U12462 ( .A(VCaptureThresh[2]), .Y(n9651) );
  INVX1 U12463 ( .A(VCaptureThresh[1]), .Y(n9648) );
  INVX1 U12464 ( .A(VCaptureThresh[0]), .Y(n9647) );
  INVX1 U12465 ( .A(ACaptureThresh[31]), .Y(n9645) );
  INVX1 U12466 ( .A(ACaptureThresh[30]), .Y(n9639) );
  INVX1 U12467 ( .A(ACaptureThresh[29]), .Y(n9637) );
  INVX1 U12468 ( .A(ACaptureThresh[28]), .Y(n9635) );
  INVX1 U12469 ( .A(ACaptureThresh[27]), .Y(n9633) );
  INVX1 U12470 ( .A(ACaptureThresh[26]), .Y(n9627) );
  INVX1 U12471 ( .A(ACaptureThresh[25]), .Y(n9625) );
  INVX1 U12472 ( .A(ACaptureThresh[24]), .Y(n9621) );
  INVX1 U12473 ( .A(ACaptureThresh[23]), .Y(n9619) );
  INVX1 U12474 ( .A(ACaptureThresh[22]), .Y(n9613) );
  INVX1 U12475 ( .A(ACaptureThresh[21]), .Y(n9611) );
  INVX1 U12476 ( .A(ACaptureThresh[20]), .Y(n9607) );
  INVX1 U12477 ( .A(ACaptureThresh[19]), .Y(n9605) );
  INVX1 U12478 ( .A(ACaptureThresh[16]), .Y(n9595) );
  INVX1 U12479 ( .A(ACaptureThresh[13]), .Y(n9585) );
  INVX1 U12480 ( .A(ACaptureThresh[12]), .Y(n9582) );
  INVX1 U12481 ( .A(ACaptureThresh[11]), .Y(n9580) );
  INVX1 U12482 ( .A(ACaptureThresh[9]), .Y(n9572) );
  INVX1 U12483 ( .A(ACaptureThresh[8]), .Y(n9567) );
  INVX1 U12484 ( .A(ACaptureThresh[7]), .Y(n9565) );
  INVX1 U12485 ( .A(ACaptureThresh[6]), .Y(n9561) );
  INVX1 U12486 ( .A(ACaptureThresh[5]), .Y(n9559) );
  INVX1 U12487 ( .A(ACaptureThresh[4]), .Y(n9557) );
  INVX1 U12488 ( .A(ACaptureThresh[3]), .Y(n9555) );
  INVX1 U12489 ( .A(ACaptureThresh[2]), .Y(n9551) );
  INVX1 U12490 ( .A(ACaptureThresh[1]), .Y(n9549) );
  INVX1 U12491 ( .A(ACaptureThresh[0]), .Y(n9548) );
  INVX1 U12492 ( .A(vflip[5]), .Y(n9545) );
  INVX1 U12493 ( .A(vflip[4]), .Y(n9544) );
  INVX1 U12494 ( .A(vflip[1]), .Y(n9541) );
  INVX1 U12495 ( .A(vflip[0]), .Y(n9533) );
  INVX1 U12496 ( .A(aflip[5]), .Y(n9493) );
  INVX1 U12497 ( .A(aflip[4]), .Y(n9492) );
  INVX1 U12498 ( .A(recentdatapoints_data_addr_reg_1533[4]), .Y(n9893) );
  INVX1 U12499 ( .A(recentdatapoints_data_addr_reg_1533[1]), .Y(n9889) );
  INVX1 U12500 ( .A(recentdatapoints_data_addr_reg_1533[0]), .Y(n9887) );
  INVX1 U12501 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][15] ), .Y(n11029) );
  INVX1 U12502 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][14] ), .Y(n11028) );
  INVX1 U12503 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][13] ), .Y(n11027) );
  INVX1 U12504 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][12] ), .Y(n11026) );
  INVX1 U12505 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][7] ), .Y(n11021) );
  INVX1 U12506 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][6] ), .Y(n11020) );
  INVX1 U12507 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][5] ), .Y(n11019) );
  INVX1 U12508 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][4] ), .Y(n11018) );
  INVX1 U12509 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][3] ), .Y(n11017) );
  INVX1 U12510 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][2] ), .Y(n11016) );
  INVX1 U12511 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][1] ), .Y(n11015) );
  INVX1 U12512 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][0] ), .Y(n11014) );
  INVX1 U12513 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][15] ), .Y(n11013) );
  INVX1 U12514 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][14] ), .Y(n11012) );
  INVX1 U12515 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][13] ), .Y(n11011) );
  INVX1 U12516 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][12] ), .Y(n11010) );
  INVX1 U12517 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][7] ), .Y(n11005) );
  INVX1 U12518 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][6] ), .Y(n11004) );
  INVX1 U12519 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][5] ), .Y(n11003) );
  INVX1 U12520 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][4] ), .Y(n11002) );
  INVX1 U12521 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][3] ), .Y(n11001) );
  INVX1 U12522 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][2] ), .Y(n11000) );
  INVX1 U12523 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][1] ), .Y(n10999) );
  INVX1 U12524 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][0] ), .Y(n10998) );
  INVX1 U12525 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][15] ), .Y(n10997) );
  INVX1 U12526 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][14] ), .Y(n10996) );
  INVX1 U12527 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][13] ), .Y(n10995) );
  INVX1 U12528 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][12] ), .Y(n10994) );
  INVX1 U12529 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][7] ), .Y(n10989) );
  INVX1 U12530 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][6] ), .Y(n10988) );
  INVX1 U12531 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][5] ), .Y(n10987) );
  INVX1 U12532 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][4] ), .Y(n10986) );
  INVX1 U12533 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][3] ), .Y(n10985) );
  INVX1 U12534 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][2] ), .Y(n10984) );
  INVX1 U12535 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][1] ), .Y(n10983) );
  INVX1 U12536 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][0] ), .Y(n10982) );
  INVX1 U12537 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][15] ), .Y(n10981) );
  INVX1 U12538 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][14] ), .Y(n10980) );
  INVX1 U12539 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][13] ), .Y(n10979) );
  INVX1 U12540 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][12] ), .Y(n10978) );
  INVX1 U12541 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][7] ), .Y(n10973) );
  INVX1 U12542 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][6] ), .Y(n10972) );
  INVX1 U12543 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][5] ), .Y(n10971) );
  INVX1 U12544 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][4] ), .Y(n10970) );
  INVX1 U12545 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][3] ), .Y(n10969) );
  INVX1 U12546 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][2] ), .Y(n10968) );
  INVX1 U12547 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][1] ), .Y(n10967) );
  INVX1 U12548 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][0] ), .Y(n10966) );
  INVX1 U12549 ( .A(aflip[1]), .Y(n9791) );
  INVX1 U12550 ( .A(aflip[0]), .Y(n9790) );
  INVX1 U12551 ( .A(VCaptureThresh[31]), .Y(n9762) );
  INVX1 U12552 ( .A(VCaptureThresh[30]), .Y(n9756) );
  INVX1 U12553 ( .A(VCaptureThresh[29]), .Y(n9754) );
  INVX1 U12554 ( .A(VCaptureThresh[28]), .Y(n9752) );
  INVX1 U12555 ( .A(VCaptureThresh[27]), .Y(n9748) );
  INVX1 U12556 ( .A(VCaptureThresh[26]), .Y(n9742) );
  INVX1 U12557 ( .A(VCaptureThresh[25]), .Y(n9739) );
  INVX1 U12558 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][11] ), .Y(n11025) );
  INVX1 U12559 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][10] ), .Y(n11024) );
  INVX1 U12560 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][9] ), .Y(n11023) );
  INVX1 U12561 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[15][8] ), .Y(n11022) );
  INVX1 U12562 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][11] ), .Y(n11009) );
  INVX1 U12563 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][10] ), .Y(n11008) );
  INVX1 U12564 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][9] ), .Y(n11007) );
  INVX1 U12565 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[7][8] ), .Y(n11006) );
  INVX1 U12566 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][11] ), .Y(n10993) );
  INVX1 U12567 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][10] ), .Y(n10992) );
  INVX1 U12568 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][9] ), .Y(n10991) );
  INVX1 U12569 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[6][8] ), .Y(n10990) );
  INVX1 U12570 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][11] ), .Y(n10977) );
  INVX1 U12571 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][10] ), .Y(n10976) );
  INVX1 U12572 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][9] ), .Y(n10975) );
  INVX1 U12573 ( .A(
        \recentdatapoints_data_U/Decision_recentdatapoints_data_ram_U/ram[4][8] ), .Y(n10974) );
  INVX1 U12574 ( .A(ACaptureThresh[18]), .Y(n9599) );
  INVX1 U12575 ( .A(ACaptureThresh[17]), .Y(n9597) );
  INVX1 U12576 ( .A(ACaptureThresh[15]), .Y(n9593) );
  INVX1 U12577 ( .A(ACaptureThresh[14]), .Y(n9587) );
  INVX1 U12578 ( .A(ACaptureThresh[10]), .Y(n9574) );
  INVX1 U12579 ( .A(CircularBuffer_len_write_assig_reg_1634[22]), .Y(n10161)
         );
  INVX1 U12580 ( .A(CircularBuffer_len_write_assig_reg_1634[21]), .Y(n10160)
         );
  INVX1 U12581 ( .A(CircularBuffer_len_write_assig_reg_1634[19]), .Y(n10158)
         );
  INVX1 U12582 ( .A(CircularBuffer_len_write_assig_reg_1634[18]), .Y(n10157)
         );
  INVX1 U12583 ( .A(CircularBuffer_len_write_assig_reg_1634[13]), .Y(n10152)
         );
  INVX1 U12584 ( .A(CircularBuffer_len_write_assig_reg_1634[12]), .Y(n10151)
         );
  INVX1 U12585 ( .A(CircularBuffer_len_write_assig_reg_1634[11]), .Y(n10150)
         );
  INVX1 U12586 ( .A(CircularBuffer_len_write_assig_reg_1634[10]), .Y(n10149)
         );
  INVX1 U12587 ( .A(CircularBuffer_len_write_assig_reg_1634[6]), .Y(n10145) );
  INVX1 U12588 ( .A(CircularBuffer_len_write_assig_2_reg_1729[22]), .Y(n10656)
         );
  INVX1 U12589 ( .A(CircularBuffer_len_write_assig_2_reg_1729[21]), .Y(n10655)
         );
  INVX1 U12590 ( .A(CircularBuffer_len_write_assig_2_reg_1729[19]), .Y(n10653)
         );
  INVX1 U12591 ( .A(CircularBuffer_len_write_assig_2_reg_1729[18]), .Y(n10652)
         );
  INVX1 U12592 ( .A(CircularBuffer_len_write_assig_2_reg_1729[13]), .Y(n10647)
         );
  INVX1 U12593 ( .A(CircularBuffer_len_write_assig_2_reg_1729[12]), .Y(n10646)
         );
  INVX1 U12594 ( .A(CircularBuffer_len_write_assig_2_reg_1729[11]), .Y(n10645)
         );
  INVX1 U12595 ( .A(CircularBuffer_len_write_assig_2_reg_1729[10]), .Y(n10644)
         );
  INVX1 U12596 ( .A(CircularBuffer_len_write_assig_2_reg_1729[6]), .Y(n10640)
         );
  INVX1 U12597 ( .A(CircularBuffer_len_read_assign_1_reg_1616[14]), .Y(n10092)
         );
  AND2X1 U12598 ( .A(s_axi_AXILiteS_AWREADY), .B(s_axi_AXILiteS_AWVALID), .Y(
        n8652) );
  INVX1 U12599 ( .A(AbeatDelay[0]), .Y(n10671) );
  INVX1 U12600 ( .A(CircularBuffer_len_read_assign_1_reg_1616[13]), .Y(n10091)
         );
  INVX1 U12601 ( .A(CircularBuffer_len_read_assign_1_reg_1616[10]), .Y(n10088)
         );
  INVX1 U12602 ( .A(CircularBuffer_len_read_assign_1_reg_1616[9]), .Y(n10087)
         );
  INVX1 U12603 ( .A(VbeatDelay[0]), .Y(n10452) );
  INVX1 U12604 ( .A(VbeatFallDelay[0]), .Y(n10365) );
  INVX1 U12605 ( .A(CircularBuffer_len_read_assign_1_reg_1616[29]), .Y(n10107)
         );
  INVX1 U12606 ( .A(CircularBuffer_len_read_assign_1_reg_1616[28]), .Y(n10106)
         );
  INVX1 U12607 ( .A(CircularBuffer_len_read_assign_1_reg_1616[25]), .Y(n10103)
         );
  INVX1 U12608 ( .A(CircularBuffer_len_read_assign_1_reg_1616[24]), .Y(n10102)
         );
  INVX1 U12609 ( .A(CircularBuffer_len_read_assign_1_reg_1616[23]), .Y(n10101)
         );
  INVX1 U12610 ( .A(CircularBuffer_len_read_assign_1_reg_1616[22]), .Y(n10100)
         );
  INVX1 U12611 ( .A(CircularBuffer_len_read_assign_1_reg_1616[8]), .Y(n10086)
         );
  INVX1 U12612 ( .A(\tmp_8_reg_1630[0] ), .Y(n10077) );
  INVX1 U12613 ( .A(recentVBools_head_i[1]), .Y(n10054) );
  INVX1 U12614 ( .A(recentVBools_head_i[2]), .Y(n10052) );
  INVX1 U12615 ( .A(recentVBools_head_i[4]), .Y(n10050) );
  INVX1 U12616 ( .A(recentVBools_head_i[3]), .Y(n9963) );
  INVX1 U12617 ( .A(CircularBuffer_len_write_assig_reg_1634[30]), .Y(n10169)
         );
  INVX1 U12618 ( .A(CircularBuffer_len_write_assig_reg_1634[29]), .Y(n10168)
         );
  INVX1 U12619 ( .A(CircularBuffer_len_write_assig_reg_1634[26]), .Y(n10165)
         );
  INVX1 U12620 ( .A(CircularBuffer_len_write_assig_reg_1634[25]), .Y(n10164)
         );
  INVX1 U12621 ( .A(CircularBuffer_len_write_assig_2_reg_1729[30]), .Y(n10664)
         );
  INVX1 U12622 ( .A(CircularBuffer_len_write_assig_2_reg_1729[29]), .Y(n10663)
         );
  INVX1 U12623 ( .A(CircularBuffer_len_write_assig_2_reg_1729[26]), .Y(n10660)
         );
  INVX1 U12624 ( .A(CircularBuffer_len_write_assig_2_reg_1729[25]), .Y(n10659)
         );
  INVX1 U12625 ( .A(n7834), .Y(n10688) );
  INVX1 U12626 ( .A(n11078), .Y(n10675) );
  INVX1 U12627 ( .A(n11079), .Y(n10685) );
  INVX1 U12628 ( .A(\Decision_AXILiteS_s_axi_U/n604 ), .Y(n9277) );
  INVX1 U12629 ( .A(tmp_38_i_reg_1550[10]), .Y(n9922) );
  INVX1 U12630 ( .A(tmp_38_i_reg_1550[22]), .Y(n9910) );
  INVX1 U12631 ( .A(tmp_38_i_reg_1550[25]), .Y(n9907) );
  INVX1 U12632 ( .A(p_tmp_i_reg_1556[4]), .Y(n9896) );
  INVX1 U12633 ( .A(recentdatapoints_head_i[2]), .Y(n9894) );
  INVX1 U12634 ( .A(recentdatapoints_head_i[4]), .Y(n9892) );
  INVX1 U12635 ( .A(recentdatapoints_head_i[3]), .Y(n9890) );
  INVX1 U12636 ( .A(recentdatapoints_head_i[1]), .Y(n9888) );
  INVX1 U12637 ( .A(recentdatapoints_len[27]), .Y(n9854) );
  INVX1 U12638 ( .A(recentdatapoints_len[26]), .Y(n9853) );
  INVX1 U12639 ( .A(recentdatapoints_len[23]), .Y(n9850) );
  INVX1 U12640 ( .A(recentdatapoints_len[22]), .Y(n9849) );
  INVX1 U12641 ( .A(recentdatapoints_len[19]), .Y(n9846) );
  INVX1 U12642 ( .A(recentdatapoints_len[16]), .Y(n9843) );
  INVX1 U12643 ( .A(recentdatapoints_len[15]), .Y(n9842) );
  INVX1 U12644 ( .A(recentdatapoints_len[9]), .Y(n9837) );
  INVX1 U12645 ( .A(recentdatapoints_len[8]), .Y(n9836) );
  INVX1 U12646 ( .A(recentdatapoints_len[4]), .Y(n9832) );
  INVX1 U12647 ( .A(recentdatapoints_len[2]), .Y(n9829) );
  INVX1 U12648 ( .A(recentdatapoints_len[1]), .Y(n9827) );
  INVX1 U12649 ( .A(recentdatapoints_len[10]), .Y(n9826) );
  OR2X1 U12650 ( .A(n9705), .B(tmp_7_reg_1544[16]), .Y(n12049) );
  INVX1 U12651 ( .A(n12025), .Y(n9670) );
  OR2X1 U12652 ( .A(n9596), .B(tmp_6_reg_1538[16]), .Y(n11960) );
  INVX1 U12653 ( .A(n11936), .Y(n9570) );
  OR2X1 U12654 ( .A(n10409), .B(VbeatDelay_new_1_reg_326[16]), .Y(n11852) );
  INVX1 U12655 ( .A(n11828), .Y(n10386) );
  OR2X1 U12656 ( .A(n10711), .B(VbeatDelay_new_1_reg_326[16]), .Y(n11128) );
  INVX1 U12657 ( .A(n11104), .Y(n10470) );
  AND2X1 U12658 ( .A(n11052), .B(n11051), .Y(n11053) );
  AND2X1 U12659 ( .A(n11072), .B(n11071), .Y(n11073) );
  INVX1 U12660 ( .A(n8066), .Y(n10398) );
  INVX1 U12661 ( .A(n8307), .Y(n10482) );
  INVX1 U12662 ( .A(n8067), .Y(n9353) );
  INVX1 U12663 ( .A(n8065), .Y(n9689) );
  INVX1 U12664 ( .A(n8064), .Y(n9583) );
  INVX1 U12665 ( .A(n7629), .Y(n9476) );
  INVX1 U12666 ( .A(n8068), .Y(n9511) );
  INVX1 U12667 ( .A(data_read_reg_1495[15]), .Y(n9793) );
  INVX1 U12668 ( .A(data_read_reg_1495[14]), .Y(n9794) );
  INVX1 U12669 ( .A(data_read_reg_1495[13]), .Y(n9795) );
  INVX1 U12670 ( .A(data_read_reg_1495[12]), .Y(n9796) );
  INVX1 U12671 ( .A(data_read_reg_1495[11]), .Y(n9797) );
  INVX1 U12672 ( .A(data_read_reg_1495[10]), .Y(n9798) );
  INVX1 U12673 ( .A(data_read_reg_1495[9]), .Y(n9799) );
  INVX1 U12674 ( .A(data_read_reg_1495[8]), .Y(n9800) );
  INVX1 U12675 ( .A(data_read_reg_1495[7]), .Y(n9801) );
  INVX1 U12676 ( .A(data_read_reg_1495[6]), .Y(n9802) );
  INVX1 U12677 ( .A(data_read_reg_1495[5]), .Y(n9803) );
  INVX1 U12678 ( .A(data_read_reg_1495[4]), .Y(n9804) );
  INVX1 U12679 ( .A(data_read_reg_1495[3]), .Y(n9805) );
  INVX1 U12680 ( .A(data_read_reg_1495[2]), .Y(n9806) );
  INVX1 U12681 ( .A(data_read_reg_1495[1]), .Y(n9807) );
  INVX1 U12682 ( .A(data_read_reg_1495[0]), .Y(n9808) );
  INVX1 U12683 ( .A(athresh[7]), .Y(n10867) );
  INVX1 U12684 ( .A(athresh[6]), .Y(n10866) );
  INVX1 U12685 ( .A(athresh[5]), .Y(n10865) );
  INVX1 U12686 ( .A(athresh[4]), .Y(n10864) );
  INVX1 U12687 ( .A(athresh[3]), .Y(n10863) );
  INVX1 U12688 ( .A(athresh[2]), .Y(n10862) );
  INVX1 U12689 ( .A(athresh[1]), .Y(n10861) );
  INVX1 U12690 ( .A(athresh[0]), .Y(n10860) );
  INVX1 U12691 ( .A(vthresh[7]), .Y(n10859) );
  INVX1 U12692 ( .A(vthresh[6]), .Y(n10858) );
  INVX1 U12693 ( .A(vthresh[5]), .Y(n10857) );
  INVX1 U12694 ( .A(vthresh[4]), .Y(n10856) );
  INVX1 U12695 ( .A(vthresh[3]), .Y(n10855) );
  INVX1 U12696 ( .A(vthresh[2]), .Y(n10854) );
  INVX1 U12697 ( .A(vthresh[1]), .Y(n10853) );
  INVX1 U12698 ( .A(vthresh[0]), .Y(n10852) );
  INVX1 U12699 ( .A(a_length[7]), .Y(n10835) );
  INVX1 U12700 ( .A(a_length[6]), .Y(n10834) );
  INVX1 U12701 ( .A(a_length[5]), .Y(n10833) );
  INVX1 U12702 ( .A(a_length[4]), .Y(n10832) );
  INVX1 U12703 ( .A(a_length[3]), .Y(n10831) );
  INVX1 U12704 ( .A(a_length[2]), .Y(n10830) );
  INVX1 U12705 ( .A(a_length[1]), .Y(n10829) );
  INVX1 U12706 ( .A(a_length[0]), .Y(n10828) );
  INVX1 U12707 ( .A(v_length[7]), .Y(n10827) );
  INVX1 U12708 ( .A(v_length[6]), .Y(n10826) );
  INVX1 U12709 ( .A(v_length[5]), .Y(n10825) );
  INVX1 U12710 ( .A(v_length[4]), .Y(n10824) );
  INVX1 U12711 ( .A(v_length[3]), .Y(n10823) );
  INVX1 U12712 ( .A(v_length[2]), .Y(n10822) );
  INVX1 U12713 ( .A(v_length[1]), .Y(n10821) );
  INVX1 U12714 ( .A(v_length[0]), .Y(n10820) );
  INVX1 U12715 ( .A(data[7]), .Y(n10819) );
  INVX1 U12716 ( .A(data[6]), .Y(n10818) );
  INVX1 U12717 ( .A(data[5]), .Y(n10817) );
  INVX1 U12718 ( .A(data[4]), .Y(n10816) );
  INVX1 U12719 ( .A(data[3]), .Y(n10815) );
  INVX1 U12720 ( .A(data[2]), .Y(n10814) );
  INVX1 U12721 ( .A(data[1]), .Y(n10813) );
  INVX1 U12722 ( .A(data[0]), .Y(n10812) );
  INVX1 U12723 ( .A(a_flip[7]), .Y(n10851) );
  INVX1 U12724 ( .A(a_flip[6]), .Y(n10850) );
  INVX1 U12725 ( .A(a_flip[5]), .Y(n10849) );
  INVX1 U12726 ( .A(a_flip[4]), .Y(n10848) );
  INVX1 U12727 ( .A(a_flip[3]), .Y(n10847) );
  INVX1 U12728 ( .A(a_flip[2]), .Y(n10846) );
  INVX1 U12729 ( .A(a_flip[1]), .Y(n10845) );
  INVX1 U12730 ( .A(a_flip[0]), .Y(n10844) );
  INVX1 U12731 ( .A(v_flip[7]), .Y(n10843) );
  INVX1 U12732 ( .A(v_flip[6]), .Y(n10842) );
  INVX1 U12733 ( .A(v_flip[5]), .Y(n10841) );
  INVX1 U12734 ( .A(v_flip[4]), .Y(n10840) );
  INVX1 U12735 ( .A(v_flip[3]), .Y(n10839) );
  INVX1 U12736 ( .A(v_flip[2]), .Y(n10838) );
  INVX1 U12737 ( .A(v_flip[1]), .Y(n10837) );
  INVX1 U12738 ( .A(v_flip[0]), .Y(n10836) );
  AND2X1 U12739 ( .A(s_axi_AXILiteS_WDATA[7]), .B(
        \Decision_AXILiteS_s_axi_U/n617 ), .Y(\Decision_AXILiteS_s_axi_U/n356 ) );
  AND2X1 U12740 ( .A(s_axi_AXILiteS_WDATA[6]), .B(
        \Decision_AXILiteS_s_axi_U/n617 ), .Y(\Decision_AXILiteS_s_axi_U/n358 ) );
  AND2X1 U12741 ( .A(s_axi_AXILiteS_WDATA[5]), .B(
        \Decision_AXILiteS_s_axi_U/n617 ), .Y(\Decision_AXILiteS_s_axi_U/n360 ) );
  AND2X1 U12742 ( .A(s_axi_AXILiteS_WDATA[4]), .B(
        \Decision_AXILiteS_s_axi_U/n617 ), .Y(\Decision_AXILiteS_s_axi_U/n362 ) );
  AND2X1 U12743 ( .A(s_axi_AXILiteS_WDATA[3]), .B(
        \Decision_AXILiteS_s_axi_U/n617 ), .Y(\Decision_AXILiteS_s_axi_U/n364 ) );
  AND2X1 U12744 ( .A(s_axi_AXILiteS_WDATA[2]), .B(
        \Decision_AXILiteS_s_axi_U/n617 ), .Y(\Decision_AXILiteS_s_axi_U/n366 ) );
  AND2X1 U12745 ( .A(s_axi_AXILiteS_WDATA[1]), .B(
        \Decision_AXILiteS_s_axi_U/n617 ), .Y(\Decision_AXILiteS_s_axi_U/n368 ) );
  INVX1 U12746 ( .A(n7841), .Y(n10273) );
  INVX1 U12747 ( .A(n7630), .Y(n9992) );
  INVX1 U12748 ( .A(\Decision_AXILiteS_s_axi_U/waddr[3] ), .Y(n10895) );
  INVX1 U12749 ( .A(recentVBools_data_addr_reg_1573[1]), .Y(n10055) );
  INVX1 U12750 ( .A(recentVBools_data_addr_reg_1573[2]), .Y(n10053) );
  INVX1 U12751 ( .A(recentVBools_data_addr_reg_1573[4]), .Y(n10051) );
  INVX1 U12752 ( .A(recentVBools_data_addr_reg_1573[0]), .Y(n10025) );
  INVX1 U12753 ( .A(recentVBools_data_addr_reg_1573[3]), .Y(n9964) );
  INVX1 U12754 ( .A(N495), .Y(n9649) );
  INVX1 U12755 ( .A(n12062), .Y(n9744) );
  INVX1 U12756 ( .A(n11973), .Y(n9631) );
  INVX1 U12757 ( .A(n11091), .Y(n10471) );
  INVX1 U12758 ( .A(n11094), .Y(n10477) );
  INVX1 U12759 ( .A(n11141), .Y(n10520) );
  INVX1 U12760 ( .A(n12012), .Y(n9671) );
  INVX1 U12761 ( .A(n12015), .Y(n9680) );
  INVX1 U12762 ( .A(n11923), .Y(n9571) );
  INVX1 U12763 ( .A(n11926), .Y(n9578) );
  INVX1 U12764 ( .A(n11815), .Y(n10387) );
  INVX1 U12765 ( .A(n11818), .Y(n10393) );
  INVX1 U12766 ( .A(n11865), .Y(n10436) );
  INVX1 U12767 ( .A(VbeatDelay_new_1_reg_326[8]), .Y(n10472) );
  AND2X1 U12768 ( .A(VstimDelay[30]), .B(n8897), .Y(\dp_cluster_0/N984 ) );
  AND2X1 U12769 ( .A(AstimDelay[30]), .B(n8898), .Y(\dp_cluster_1/N952 ) );
  INVX1 U12770 ( .A(AbeatDelay_new_reg_394[31]), .Y(n10741) );
  BUFX2 U12771 ( .A(s_axi_AXILiteS_ARADDR[5]), .Y(n8859) );
  INVX1 U12772 ( .A(a_thresh[29]), .Y(n9789) );
  INVX1 U12773 ( .A(a_thresh[28]), .Y(n9788) );
  INVX1 U12774 ( .A(v_thresh[29]), .Y(n9531) );
  INVX1 U12775 ( .A(v_thresh[28]), .Y(n9530) );
  AND2X1 U12776 ( .A(ap_CS_fsm[13]), .B(n5949), .Y(n8653) );
  INVX1 U12777 ( .A(CircularBuffer_len_read_assign_3_reg_1711[2]), .Y(n10575)
         );
  INVX1 U12778 ( .A(CircularBuffer_len_read_assign_1_reg_1616[2]), .Y(n10080)
         );
  INVX1 U12779 ( .A(CircularBuffer_len_read_assign_3_reg_1711[4]), .Y(n10577)
         );
  INVX1 U12780 ( .A(CircularBuffer_len_read_assign_1_reg_1616[4]), .Y(n10082)
         );
  AND2X1 U12781 ( .A(ap_CS_fsm[13]), .B(n5950), .Y(n8654) );
  INVX1 U12782 ( .A(CircularBuffer_len_read_assign_3_reg_1711[3]), .Y(n10576)
         );
  INVX1 U12783 ( .A(CircularBuffer_len_read_assign_1_reg_1616[3]), .Y(n10081)
         );
  INVX1 U12784 ( .A(ACaptureThresh_loc_reg_288[6]), .Y(n9564) );
  INVX1 U12785 ( .A(VCaptureThresh_loc_reg_298[22]), .Y(n9730) );
  INVX1 U12786 ( .A(ACaptureThresh_loc_reg_288[18]), .Y(n9604) );
  INVX1 U12787 ( .A(ACaptureThresh_loc_reg_288[22]), .Y(n9618) );
  INVX1 U12788 ( .A(VCaptureThresh_loc_reg_298[6]), .Y(n9665) );
  INVX1 U12789 ( .A(VCaptureThresh_loc_reg_298[18]), .Y(n9713) );
  INVX1 U12790 ( .A(s_axi_AXILiteS_WVALID), .Y(n9280) );
  BUFX2 U12791 ( .A(s_axi_AXILiteS_ARADDR[3]), .Y(n8858) );
  INVX1 U12792 ( .A(CircularBuffer_len_read_assign_3_reg_1711[31]), .Y(n10604)
         );
  INVX1 U12793 ( .A(CircularBuffer_len_read_assign_1_reg_1616[31]), .Y(n10109)
         );
  INVX1 U12794 ( .A(ACaptureThresh_loc_reg_288[30]), .Y(n9644) );
  INVX1 U12795 ( .A(ACaptureThresh_loc_reg_288[14]), .Y(n9592) );
  INVX1 U12796 ( .A(VCaptureThresh_loc_reg_298[14]), .Y(n9699) );
  INVX1 U12797 ( .A(ACaptureThresh_loc_reg_288[26]), .Y(n9632) );
  INVX1 U12798 ( .A(VCaptureThresh_loc_reg_298[30]), .Y(n9761) );
  INVX1 U12799 ( .A(VCaptureThresh_loc_reg_298[26]), .Y(n9747) );
  AND2X1 U12800 ( .A(\reset_params_V[0] ), .B(n8967), .Y(n8655) );
  INVX1 U12801 ( .A(ACaptureThresh_loc_reg_288[10]), .Y(n9579) );
  INVX1 U12802 ( .A(VCaptureThresh_loc_reg_298[10]), .Y(n9683) );
  AND2X1 U12803 ( .A(\tmp_8_reg_1630[0] ), .B(n9012), .Y(n8656) );
  AND2X1 U12804 ( .A(\tmp_13_reg_1725[0] ), .B(ap_CS_fsm[12]), .Y(n8657) );
  INVX1 U12805 ( .A(VbeatDelay_new_1_reg_326[7]), .Y(n10468) );
  INVX1 U12806 ( .A(ACaptureThresh_loc_reg_288[31]), .Y(n9646) );
  INVX1 U12807 ( .A(VCaptureThresh_loc_reg_298[31]), .Y(n9765) );
  AND2X1 U12808 ( .A(ap_start), .B(ap_CS_fsm[0]), .Y(n8658) );
  INVX1 U12809 ( .A(CircularBuffer_len_write_assig_2_reg_1729[1]), .Y(n10635)
         );
  INVX1 U12810 ( .A(CircularBuffer_len_write_assig_reg_1634[1]), .Y(n10140) );
  INVX1 U12811 ( .A(sum_phi_fu_311_p4[1]), .Y(n10061) );
  INVX1 U12812 ( .A(\Decision_AXILiteS_s_axi_U/n323 ), .Y(n9318) );
  INVX1 U12813 ( .A(\Decision_AXILiteS_s_axi_U/n325 ), .Y(n9313) );
  INVX1 U12814 ( .A(ap_CS_fsm[2]), .Y(n9933) );
  INVX1 U12815 ( .A(VCaptureThresh_loc_reg_298[5]), .Y(n9661) );
  INVX1 U12816 ( .A(ACaptureThresh_loc_reg_288[5]), .Y(n9560) );
  INVX1 U12817 ( .A(CircularBuffer_len_write_assig_2_reg_1729[3]), .Y(n10637)
         );
  INVX1 U12818 ( .A(CircularBuffer_len_write_assig_reg_1634[3]), .Y(n10142) );
  INVX1 U12819 ( .A(\Decision_AXILiteS_s_axi_U/n338 ), .Y(n9312) );
  INVX1 U12820 ( .A(CircularBuffer_len_write_assig_2_reg_1729[4]), .Y(n10638)
         );
  INVX1 U12821 ( .A(CircularBuffer_len_write_assig_reg_1634[4]), .Y(n10143) );
  INVX1 U12822 ( .A(ACaptureThresh_loc_reg_288[2]), .Y(n9554) );
  INVX1 U12823 ( .A(VCaptureThresh_loc_reg_298[2]), .Y(n9654) );
  INVX1 U12824 ( .A(VbeatDelay_new_1_reg_326[19]), .Y(n10501) );
  INVX1 U12825 ( .A(VbeatDelay_new_1_reg_326[15]), .Y(n10491) );
  INVX1 U12826 ( .A(\Decision_AXILiteS_s_axi_U/waddr[4] ), .Y(n10897) );
  INVX1 U12827 ( .A(p_tmp_i_reg_1556[0]), .Y(n9900) );
  AND2X1 U12828 ( .A(s_axi_AXILiteS_WSTRB[1]), .B(ap_rst_n), .Y(
        \Decision_AXILiteS_s_axi_U/n353 ) );
  INVX1 U12829 ( .A(VCaptureThresh_loc_reg_298[17]), .Y(n9707) );
  INVX1 U12830 ( .A(VCaptureThresh_loc_reg_298[21]), .Y(n9724) );
  INVX1 U12831 ( .A(ACaptureThresh_loc_reg_288[17]), .Y(n9598) );
  INVX1 U12832 ( .A(ACaptureThresh_loc_reg_288[21]), .Y(n9612) );
  INVX1 U12833 ( .A(n11262), .Y(n10302) );
  INVX1 U12834 ( .A(n11366), .Y(n10020) );
  INVX1 U12835 ( .A(n11418), .Y(n10329) );
  INVX1 U12836 ( .A(n11314), .Y(n9988) );
  INVX1 U12837 ( .A(n11266), .Y(n10300) );
  INVX1 U12838 ( .A(n11370), .Y(n10018) );
  INVX1 U12839 ( .A(n11422), .Y(n10327) );
  INVX1 U12840 ( .A(n11318), .Y(n9986) );
  INVX1 U12841 ( .A(n11270), .Y(n10298) );
  INVX1 U12842 ( .A(n11374), .Y(n10016) );
  INVX1 U12843 ( .A(n11426), .Y(n10325) );
  INVX1 U12844 ( .A(n11322), .Y(n9984) );
  INVX1 U12845 ( .A(n11274), .Y(n10296) );
  INVX1 U12846 ( .A(n11378), .Y(n10014) );
  INVX1 U12847 ( .A(n11430), .Y(n10323) );
  INVX1 U12848 ( .A(n11326), .Y(n9982) );
  INVX1 U12849 ( .A(n11278), .Y(n10294) );
  INVX1 U12850 ( .A(n11382), .Y(n10012) );
  INVX1 U12851 ( .A(n11434), .Y(n10321) );
  INVX1 U12852 ( .A(n11330), .Y(n9980) );
  INVX1 U12853 ( .A(n11282), .Y(n10292) );
  INVX1 U12854 ( .A(n11386), .Y(n10010) );
  INVX1 U12855 ( .A(n11438), .Y(n10319) );
  INVX1 U12856 ( .A(n11334), .Y(n9978) );
  INVX1 U12857 ( .A(n11286), .Y(n10290) );
  INVX1 U12858 ( .A(n11390), .Y(n10008) );
  INVX1 U12859 ( .A(n11442), .Y(n10317) );
  INVX1 U12860 ( .A(n11338), .Y(n9976) );
  INVX1 U12861 ( .A(n11290), .Y(n10288) );
  INVX1 U12862 ( .A(n11394), .Y(n10006) );
  INVX1 U12863 ( .A(n11446), .Y(n10315) );
  INVX1 U12864 ( .A(n11342), .Y(n9974) );
  INVX1 U12865 ( .A(n11294), .Y(n10286) );
  INVX1 U12866 ( .A(n11398), .Y(n10004) );
  INVX1 U12867 ( .A(n11450), .Y(n10313) );
  INVX1 U12868 ( .A(n11346), .Y(n9972) );
  INVX1 U12869 ( .A(n11298), .Y(n10284) );
  INVX1 U12870 ( .A(n11402), .Y(n10002) );
  INVX1 U12871 ( .A(n11454), .Y(n10311) );
  INVX1 U12872 ( .A(n11350), .Y(n9970) );
  INVX1 U12873 ( .A(n11302), .Y(n10282) );
  INVX1 U12874 ( .A(n11406), .Y(n10000) );
  INVX1 U12875 ( .A(n11458), .Y(n10309) );
  INVX1 U12876 ( .A(n11354), .Y(n9968) );
  INVX1 U12877 ( .A(VCaptureThresh_loc_reg_298[25]), .Y(n9741) );
  INVX1 U12878 ( .A(ACaptureThresh_loc_reg_288[25]), .Y(n9626) );
  AND2X1 U12879 ( .A(n8897), .B(VstimDelay[9]), .Y(\dp_cluster_0/N963 ) );
  AND2X1 U12880 ( .A(n8898), .B(AstimDelay[9]), .Y(\dp_cluster_1/N931 ) );
  AND2X1 U12881 ( .A(VstimDelay[1]), .B(n8897), .Y(\dp_cluster_0/N955 ) );
  AND2X1 U12882 ( .A(AstimDelay[1]), .B(n8898), .Y(\dp_cluster_1/N923 ) );
  AND2X1 U12883 ( .A(VstimDelay[2]), .B(n8897), .Y(\dp_cluster_0/N956 ) );
  AND2X1 U12884 ( .A(AstimDelay[2]), .B(n8898), .Y(\dp_cluster_1/N924 ) );
  AND2X1 U12885 ( .A(VstimDelay[3]), .B(n8897), .Y(\dp_cluster_0/N957 ) );
  AND2X1 U12886 ( .A(AstimDelay[3]), .B(n8898), .Y(\dp_cluster_1/N925 ) );
  AND2X1 U12887 ( .A(VstimDelay[4]), .B(n8897), .Y(\dp_cluster_0/N958 ) );
  AND2X1 U12888 ( .A(AstimDelay[4]), .B(n8898), .Y(\dp_cluster_1/N926 ) );
  AND2X1 U12889 ( .A(VstimDelay[5]), .B(n8897), .Y(\dp_cluster_0/N959 ) );
  AND2X1 U12890 ( .A(AstimDelay[5]), .B(n8898), .Y(\dp_cluster_1/N927 ) );
  AND2X1 U12891 ( .A(VstimDelay[6]), .B(n8897), .Y(\dp_cluster_0/N960 ) );
  AND2X1 U12892 ( .A(AstimDelay[6]), .B(n8898), .Y(\dp_cluster_1/N928 ) );
  AND2X1 U12893 ( .A(VstimDelay[7]), .B(n8897), .Y(\dp_cluster_0/N961 ) );
  AND2X1 U12894 ( .A(AstimDelay[7]), .B(n8898), .Y(\dp_cluster_1/N929 ) );
  AND2X1 U12895 ( .A(VstimDelay[8]), .B(n8897), .Y(\dp_cluster_0/N962 ) );
  AND2X1 U12896 ( .A(AstimDelay[8]), .B(n8898), .Y(\dp_cluster_1/N930 ) );
  AND2X1 U12897 ( .A(VstimDelay[10]), .B(n8897), .Y(\dp_cluster_0/N964 ) );
  AND2X1 U12898 ( .A(AstimDelay[10]), .B(n8898), .Y(\dp_cluster_1/N932 ) );
  AND2X1 U12899 ( .A(VstimDelay[11]), .B(n8897), .Y(\dp_cluster_0/N965 ) );
  AND2X1 U12900 ( .A(AstimDelay[11]), .B(n8898), .Y(\dp_cluster_1/N933 ) );
  AND2X1 U12901 ( .A(VstimDelay[12]), .B(n8897), .Y(\dp_cluster_0/N966 ) );
  AND2X1 U12902 ( .A(AstimDelay[12]), .B(n8898), .Y(\dp_cluster_1/N934 ) );
  AND2X1 U12903 ( .A(VstimDelay[13]), .B(n8897), .Y(\dp_cluster_0/N967 ) );
  AND2X1 U12904 ( .A(AstimDelay[13]), .B(n8898), .Y(\dp_cluster_1/N935 ) );
  AND2X1 U12905 ( .A(VstimDelay[14]), .B(n8897), .Y(\dp_cluster_0/N968 ) );
  AND2X1 U12906 ( .A(AstimDelay[14]), .B(n8898), .Y(\dp_cluster_1/N936 ) );
  AND2X1 U12907 ( .A(VstimDelay[15]), .B(n8897), .Y(\dp_cluster_0/N969 ) );
  AND2X1 U12908 ( .A(AstimDelay[15]), .B(n8898), .Y(\dp_cluster_1/N937 ) );
  AND2X1 U12909 ( .A(VstimDelay[16]), .B(n8897), .Y(\dp_cluster_0/N970 ) );
  AND2X1 U12910 ( .A(AstimDelay[16]), .B(n8898), .Y(\dp_cluster_1/N938 ) );
  AND2X1 U12911 ( .A(VstimDelay[17]), .B(n8897), .Y(\dp_cluster_0/N971 ) );
  AND2X1 U12912 ( .A(AstimDelay[17]), .B(n8898), .Y(\dp_cluster_1/N939 ) );
  AND2X1 U12913 ( .A(VstimDelay[18]), .B(n8897), .Y(\dp_cluster_0/N972 ) );
  AND2X1 U12914 ( .A(AstimDelay[18]), .B(n8898), .Y(\dp_cluster_1/N940 ) );
  AND2X1 U12915 ( .A(VstimDelay[19]), .B(n8897), .Y(\dp_cluster_0/N973 ) );
  AND2X1 U12916 ( .A(AstimDelay[19]), .B(n8898), .Y(\dp_cluster_1/N941 ) );
  AND2X1 U12917 ( .A(VstimDelay[20]), .B(n8897), .Y(\dp_cluster_0/N974 ) );
  AND2X1 U12918 ( .A(AstimDelay[20]), .B(n8898), .Y(\dp_cluster_1/N942 ) );
  AND2X1 U12919 ( .A(VstimDelay[21]), .B(n8897), .Y(\dp_cluster_0/N975 ) );
  AND2X1 U12920 ( .A(AstimDelay[21]), .B(n8898), .Y(\dp_cluster_1/N943 ) );
  AND2X1 U12921 ( .A(VstimDelay[22]), .B(n8897), .Y(\dp_cluster_0/N976 ) );
  AND2X1 U12922 ( .A(AstimDelay[22]), .B(n8898), .Y(\dp_cluster_1/N944 ) );
  AND2X1 U12923 ( .A(VstimDelay[23]), .B(n8897), .Y(\dp_cluster_0/N977 ) );
  AND2X1 U12924 ( .A(AstimDelay[23]), .B(n8898), .Y(\dp_cluster_1/N945 ) );
  AND2X1 U12925 ( .A(VstimDelay[24]), .B(n8897), .Y(\dp_cluster_0/N978 ) );
  AND2X1 U12926 ( .A(AstimDelay[24]), .B(n8898), .Y(\dp_cluster_1/N946 ) );
  AND2X1 U12927 ( .A(VstimDelay[25]), .B(n8897), .Y(\dp_cluster_0/N979 ) );
  AND2X1 U12928 ( .A(AstimDelay[25]), .B(n8898), .Y(\dp_cluster_1/N947 ) );
  AND2X1 U12929 ( .A(VstimDelay[26]), .B(n8897), .Y(\dp_cluster_0/N980 ) );
  AND2X1 U12930 ( .A(AstimDelay[26]), .B(n8898), .Y(\dp_cluster_1/N948 ) );
  AND2X1 U12931 ( .A(VstimDelay[27]), .B(n8897), .Y(\dp_cluster_0/N981 ) );
  AND2X1 U12932 ( .A(AstimDelay[27]), .B(n8898), .Y(\dp_cluster_1/N949 ) );
  AND2X1 U12933 ( .A(VstimDelay[28]), .B(n8897), .Y(\dp_cluster_0/N982 ) );
  AND2X1 U12934 ( .A(AstimDelay[28]), .B(n8898), .Y(\dp_cluster_1/N950 ) );
  AND2X1 U12935 ( .A(VstimDelay[29]), .B(n8897), .Y(\dp_cluster_0/N983 ) );
  AND2X1 U12936 ( .A(AstimDelay[29]), .B(n8898), .Y(\dp_cluster_1/N951 ) );
  INVX1 U12937 ( .A(VCaptureThresh_loc_reg_298[13]), .Y(n9693) );
  INVX1 U12938 ( .A(VCaptureThresh_loc_reg_298[29]), .Y(n9755) );
  INVX1 U12939 ( .A(ACaptureThresh_loc_reg_288[13]), .Y(n9586) );
  INVX1 U12940 ( .A(ACaptureThresh_loc_reg_288[29]), .Y(n9638) );
  BUFX2 U12941 ( .A(s_axi_AXILiteS_ARADDR[2]), .Y(n8857) );
  INVX1 U12942 ( .A(CircularBuffer_len_write_assig_2_reg_1729[31]), .Y(n10665)
         );
  INVX1 U12943 ( .A(CircularBuffer_len_write_assig_reg_1634[31]), .Y(n10170)
         );
  INVX1 U12944 ( .A(VbeatDelay_new_1_reg_326[27]), .Y(n10523) );
  INVX1 U12945 ( .A(VbeatDelay_new_1_reg_326[23]), .Y(n10512) );
  INVX1 U12946 ( .A(CircularBuffer_len_write_assig_2_reg_1729[2]), .Y(n10636)
         );
  INVX1 U12947 ( .A(CircularBuffer_len_write_assig_reg_1634[2]), .Y(n10141) );
  INVX1 U12948 ( .A(VbeatDelay_new_1_reg_326[3]), .Y(n10459) );
  INVX1 U12949 ( .A(VbeatDelay_new_1_reg_326[11]), .Y(n10480) );
  OR2X1 U12950 ( .A(n9042), .B(s_axi_AXILiteS_WSTRB[1]), .Y(
        \Decision_AXILiteS_s_axi_U/n352 ) );
  INVX1 U12951 ( .A(\Decision_AXILiteS_s_axi_U/waddr[6] ), .Y(n10899) );
  INVX1 U12952 ( .A(\Decision_AXILiteS_s_axi_U/waddr[5] ), .Y(n10898) );
  INVX1 U12953 ( .A(s_axi_AXILiteS_WDATA[15]), .Y(n9298) );
  INVX1 U12954 ( .A(s_axi_AXILiteS_WDATA[14]), .Y(n9299) );
  INVX1 U12955 ( .A(s_axi_AXILiteS_WDATA[13]), .Y(n9300) );
  INVX1 U12956 ( .A(s_axi_AXILiteS_WDATA[12]), .Y(n9301) );
  INVX1 U12957 ( .A(s_axi_AXILiteS_WDATA[11]), .Y(n9302) );
  INVX1 U12958 ( .A(s_axi_AXILiteS_WDATA[10]), .Y(n9303) );
  INVX1 U12959 ( .A(s_axi_AXILiteS_WDATA[9]), .Y(n9304) );
  INVX1 U12960 ( .A(s_axi_AXILiteS_WDATA[8]), .Y(n9305) );
  INVX1 U12961 ( .A(AbeatDelay_new_reg_394[22]), .Y(n10723) );
  INVX1 U12962 ( .A(s_axi_AXILiteS_ARADDR[4]), .Y(n9319) );
  AND2X1 U12963 ( .A(s_axi_AXILiteS_WSTRB[2]), .B(ap_rst_n), .Y(
        \Decision_AXILiteS_s_axi_U/n397 ) );
  INVX1 U12964 ( .A(ACaptureThresh_loc_reg_288[24]), .Y(n9624) );
  INVX1 U12965 ( .A(VCaptureThresh_loc_reg_298[24]), .Y(n9738) );
  INVX1 U12966 ( .A(AbeatDelay_new_reg_394[30]), .Y(n10739) );
  AND2X1 U12967 ( .A(s_axi_AXILiteS_WSTRB[3]), .B(ap_rst_n), .Y(
        \Decision_AXILiteS_s_axi_U/n385 ) );
  INVX1 U12968 ( .A(AbeatDelay_new_reg_394[18]), .Y(n10715) );
  INVX1 U12969 ( .A(AbeatDelay_new_reg_394[2]), .Y(n10681) );
  INVX1 U12970 ( .A(CircularBuffer_len_write_assig_3_fu_1249_p2[0]), .Y(n10541) );
  INVX1 U12971 ( .A(CircularBuffer_len_write_assig_1_fu_924_p2[0]), .Y(n10076)
         );
  INVX1 U12972 ( .A(AbeatDelay_new_reg_394[6]), .Y(n10691) );
  INVX1 U12973 ( .A(AbeatDelay_new_reg_394[7]), .Y(n10693) );
  INVX1 U12974 ( .A(CircularBuffer_len_read_assign_3_reg_1711[5]), .Y(n10578)
         );
  INVX1 U12975 ( .A(CircularBuffer_len_read_assign_1_reg_1616[5]), .Y(n10083)
         );
  INVX1 U12976 ( .A(CircularBuffer_len_write_assig_2_reg_1729[0]), .Y(n10634)
         );
  INVX1 U12977 ( .A(CircularBuffer_len_write_assig_reg_1634[0]), .Y(n10139) );
  INVX1 U12978 ( .A(VbeatFallDelay_new_1_reg_342[31]), .Y(n10449) );
  INVX1 U12979 ( .A(AbeatDelay_new_reg_394[26]), .Y(n10731) );
  INVX1 U12980 ( .A(AbeatDelay_new_reg_394[14]), .Y(n10707) );
  INVX1 U12981 ( .A(AbeatDelay_new_reg_394[10]), .Y(n10699) );
  INVX1 U12982 ( .A(AbeatDelay_new_reg_394[17]), .Y(n10713) );
  INVX1 U12983 ( .A(AbeatDelay_new_reg_394[21]), .Y(n10721) );
  INVX1 U12984 ( .A(AbeatDelay_new_reg_394[20]), .Y(n10719) );
  INVX1 U12985 ( .A(AbeatDelay_new_reg_394[5]), .Y(n10689) );
  INVX1 U12986 ( .A(VCaptureThresh_loc_reg_298[12]), .Y(n9690) );
  INVX1 U12987 ( .A(VCaptureThresh_loc_reg_298[28]), .Y(n9753) );
  INVX1 U12988 ( .A(ACaptureThresh_loc_reg_288[12]), .Y(n9584) );
  INVX1 U12989 ( .A(ACaptureThresh_loc_reg_288[28]), .Y(n9636) );
  INVX1 U12990 ( .A(AbeatDelay_new_reg_394[1]), .Y(n10679) );
  INVX1 U12991 ( .A(recentABools_head_i[0]), .Y(n10271) );
  XNOR2X1 U12992 ( .A(\add_1405/carry[31] ), .B(recentdatapoints_head_i[31]), 
        .Y(n8659) );
  XNOR2X1 U12993 ( .A(\add_1393/carry[31] ), .B(recentVBools_head_i[31]), .Y(
        n8660) );
  XNOR2X1 U12994 ( .A(\add_1391/carry[31] ), .B(recentABools_head_i[31]), .Y(
        n8661) );
  INVX1 U12995 ( .A(recentVBools_head_i[0]), .Y(n10024) );
  INVX1 U12996 ( .A(AbeatDelay_new_reg_394[24]), .Y(n10727) );
  INVX1 U12997 ( .A(AbeatDelay_new_reg_394[9]), .Y(n10697) );
  INVX1 U12998 ( .A(tmp_7_reg_1544[8]), .Y(n10785) );
  INVX1 U12999 ( .A(tmp_6_reg_1538[8]), .Y(n10751) );
  INVX1 U13000 ( .A(VbeatDelay_new_1_reg_326[1]), .Y(n10454) );
  INVX1 U13001 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[6]), .Y(n10333)
         );
  INVX1 U13002 ( .A(CircularBuffer_head_i_read_ass_reg_1624[6]), .Y(n10026) );
  INVX1 U13003 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[9]), .Y(n10335)
         );
  INVX1 U13004 ( .A(CircularBuffer_head_i_read_ass_reg_1624[9]), .Y(n10028) );
  INVX1 U13005 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[11]), .Y(n10337)
         );
  INVX1 U13006 ( .A(CircularBuffer_head_i_read_ass_reg_1624[11]), .Y(n10030)
         );
  INVX1 U13007 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[13]), .Y(n10339)
         );
  INVX1 U13008 ( .A(CircularBuffer_head_i_read_ass_reg_1624[13]), .Y(n10032)
         );
  INVX1 U13009 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[15]), .Y(n10341)
         );
  INVX1 U13010 ( .A(CircularBuffer_head_i_read_ass_reg_1624[15]), .Y(n10034)
         );
  INVX1 U13011 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[17]), .Y(n10343)
         );
  INVX1 U13012 ( .A(CircularBuffer_head_i_read_ass_reg_1624[17]), .Y(n10036)
         );
  INVX1 U13013 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[19]), .Y(n10345)
         );
  INVX1 U13014 ( .A(CircularBuffer_head_i_read_ass_reg_1624[19]), .Y(n10038)
         );
  INVX1 U13015 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[21]), .Y(n10347)
         );
  INVX1 U13016 ( .A(CircularBuffer_head_i_read_ass_reg_1624[21]), .Y(n10040)
         );
  INVX1 U13017 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[23]), .Y(n10349)
         );
  INVX1 U13018 ( .A(CircularBuffer_head_i_read_ass_reg_1624[23]), .Y(n10042)
         );
  INVX1 U13019 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[25]), .Y(n10351)
         );
  INVX1 U13020 ( .A(CircularBuffer_head_i_read_ass_reg_1624[25]), .Y(n10044)
         );
  INVX1 U13021 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[27]), .Y(n10353)
         );
  INVX1 U13022 ( .A(CircularBuffer_head_i_read_ass_reg_1624[27]), .Y(n10046)
         );
  INVX1 U13023 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[30]), .Y(n10356)
         );
  INVX1 U13024 ( .A(CircularBuffer_head_i_read_ass_reg_1624[30]), .Y(n10049)
         );
  INVX1 U13025 ( .A(AbeatDelay_new_reg_394[28]), .Y(n10735) );
  OR2X1 U13026 ( .A(n9042), .B(s_axi_AXILiteS_WSTRB[3]), .Y(
        \Decision_AXILiteS_s_axi_U/n384 ) );
  OR2X1 U13027 ( .A(n9042), .B(s_axi_AXILiteS_WSTRB[2]), .Y(
        \Decision_AXILiteS_s_axi_U/n396 ) );
  INVX1 U13028 ( .A(AbeatDelay_new_reg_394[16]), .Y(n10711) );
  INVX1 U13029 ( .A(VbeatDelay_new_1_reg_326[30]), .Y(n10531) );
  INVX1 U13030 ( .A(p_tmp_i_reg_1556[2]), .Y(n9898) );
  INVX1 U13031 ( .A(p_tmp_i_reg_1556[3]), .Y(n9897) );
  INVX1 U13032 ( .A(p_tmp_i_reg_1556[1]), .Y(n9899) );
  INVX1 U13033 ( .A(AbeatDelay_new_reg_394[8]), .Y(n10695) );
  INVX1 U13034 ( .A(VbeatDelay_new_1_reg_326[22]), .Y(n10510) );
  INVX1 U13035 ( .A(VbeatDelay_new_1_reg_326[6]), .Y(n10466) );
  INVX1 U13036 ( .A(VbeatDelay_new_1_reg_326[2]), .Y(n10457) );
  INVX1 U13037 ( .A(VbeatDelay_new_1_reg_326[26]), .Y(n10521) );
  INVX1 U13038 ( .A(AbeatDelay_new_reg_394[12]), .Y(n10703) );
  INVX1 U13039 ( .A(VbeatDelay_new_1_reg_326[14]), .Y(n10489) );
  INVX1 U13040 ( .A(VbeatDelay_new_1_reg_326[18]), .Y(n10499) );
  INVX1 U13041 ( .A(VCaptureThresh_loc_reg_298[4]), .Y(n9659) );
  INVX1 U13042 ( .A(ACaptureThresh_loc_reg_288[4]), .Y(n9558) );
  INVX1 U13043 ( .A(AbeatDelay_new_reg_394[4]), .Y(n10686) );
  INVX1 U13044 ( .A(VbeatFallDelay_new_1_reg_342[10]), .Y(n10394) );
  XNOR2X1 U13045 ( .A(\tmp_12_reg_1694[0] ), .B(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[0]), .Y(n8662) );
  XNOR2X1 U13046 ( .A(\tmp_s_reg_1578[0] ), .B(
        CircularBuffer_int_30_sum_i_fu_758_p3[0]), .Y(n8663) );
  INVX1 U13047 ( .A(AbeatDelay_new_reg_394[29]), .Y(n10737) );
  INVX1 U13048 ( .A(AbeatDelay_new_reg_394[25]), .Y(n10729) );
  INVX1 U13049 ( .A(AbeatDelay_new_reg_394[13]), .Y(n10705) );
  INVX1 U13050 ( .A(n11538), .Y(n9733) );
  INVX1 U13051 ( .A(ACaptureThresh_loc_reg_288[7]), .Y(n9566) );
  INVX1 U13052 ( .A(ACaptureThresh_loc_reg_288[3]), .Y(n9556) );
  INVX1 U13053 ( .A(ACaptureThresh_loc_reg_288[11]), .Y(n9581) );
  INVX1 U13054 ( .A(ACaptureThresh_loc_reg_288[15]), .Y(n9594) );
  INVX1 U13055 ( .A(ACaptureThresh_loc_reg_288[19]), .Y(n9606) );
  INVX1 U13056 ( .A(ACaptureThresh_loc_reg_288[23]), .Y(n9620) );
  INVX1 U13057 ( .A(ACaptureThresh_loc_reg_288[27]), .Y(n9634) );
  INVX1 U13058 ( .A(VCaptureThresh_loc_reg_298[7]), .Y(n9668) );
  INVX1 U13059 ( .A(VCaptureThresh_loc_reg_298[3]), .Y(n9657) );
  INVX1 U13060 ( .A(VCaptureThresh_loc_reg_298[11]), .Y(n9687) );
  INVX1 U13061 ( .A(VCaptureThresh_loc_reg_298[15]), .Y(n9703) );
  INVX1 U13062 ( .A(VCaptureThresh_loc_reg_298[19]), .Y(n9717) );
  INVX1 U13063 ( .A(VCaptureThresh_loc_reg_298[23]), .Y(n9734) );
  INVX1 U13064 ( .A(VCaptureThresh_loc_reg_298[27]), .Y(n9751) );
  INVX1 U13065 ( .A(n12007), .Y(n9695) );
  INVX1 U13066 ( .A(n12052), .Y(n9757) );
  INVX1 U13067 ( .A(n11918), .Y(n9590) );
  INVX1 U13068 ( .A(n11963), .Y(n9642) );
  INVX1 U13069 ( .A(VbeatDelay_new_1_reg_326[31]), .Y(n10533) );
  AND2X1 U13070 ( .A(AstimDelay[0]), .B(n8898), .Y(\dp_cluster_1/N922 ) );
  AND2X1 U13071 ( .A(VstimDelay[0]), .B(n8897), .Y(\dp_cluster_0/N954 ) );
  INVX1 U13072 ( .A(n11841), .Y(n10381) );
  INVX1 U13073 ( .A(VbeatDelay_new_1_reg_326[12]), .Y(n10483) );
  INVX1 U13074 ( .A(n11707), .Y(n9615) );
  INVX1 U13075 ( .A(n12171), .Y(n9729) );
  INVX1 U13076 ( .A(n12038), .Y(n9663) );
  INVX1 U13077 ( .A(n11949), .Y(n9563) );
  INVX1 U13078 ( .A(n11745), .Y(n9376) );
  INVX1 U13079 ( .A(n11487), .Y(n9656) );
  INVX1 U13080 ( .A(VCaptureThresh_loc_reg_298[9]), .Y(n9677) );
  INVX1 U13081 ( .A(ACaptureThresh_loc_reg_288[9]), .Y(n9573) );
  INVX1 U13082 ( .A(n11834), .Y(n10372) );
  INVX1 U13083 ( .A(VbeatDelay_new_1_reg_326[21]), .Y(n10506) );
  INVX1 U13084 ( .A(VbeatDelay_new_1_reg_326[5]), .Y(n10463) );
  INVX1 U13085 ( .A(n11810), .Y(n10403) );
  INVX1 U13086 ( .A(n11855), .Y(n10445) );
  INVX1 U13087 ( .A(n11086), .Y(n10487) );
  INVX1 U13088 ( .A(n11131), .Y(n10529) );
  INVX1 U13089 ( .A(n11117), .Y(n10465) );
  INVX1 U13090 ( .A(n11752), .Y(n9370) );
  INVX1 U13091 ( .A(n11656), .Y(n9552) );
  INVX1 U13092 ( .A(n12120), .Y(n9653) );
  INVX1 U13093 ( .A(n12031), .Y(n9652) );
  INVX1 U13094 ( .A(n11942), .Y(n9553) );
  INVX1 U13095 ( .A(ap_CS_fsm[5]), .Y(n10056) );
  INVX1 U13096 ( .A(tmp_7_reg_1544[7]), .Y(n10784) );
  INVX1 U13097 ( .A(tmp_7_reg_1544[3]), .Y(n10780) );
  INVX1 U13098 ( .A(tmp_7_reg_1544[11]), .Y(n10788) );
  INVX1 U13099 ( .A(tmp_7_reg_1544[15]), .Y(n10792) );
  INVX1 U13100 ( .A(tmp_7_reg_1544[27]), .Y(n10804) );
  INVX1 U13101 ( .A(tmp_6_reg_1538[7]), .Y(n10750) );
  INVX1 U13102 ( .A(tmp_6_reg_1538[3]), .Y(n10746) );
  INVX1 U13103 ( .A(tmp_6_reg_1538[11]), .Y(n10754) );
  INVX1 U13104 ( .A(tmp_6_reg_1538[15]), .Y(n10758) );
  INVX1 U13105 ( .A(tmp_6_reg_1538[27]), .Y(n10770) );
  INVX1 U13106 ( .A(tmp_7_reg_1544[19]), .Y(n10796) );
  INVX1 U13107 ( .A(tmp_7_reg_1544[23]), .Y(n10800) );
  INVX1 U13108 ( .A(tmp_6_reg_1538[19]), .Y(n10762) );
  INVX1 U13109 ( .A(tmp_6_reg_1538[23]), .Y(n10766) );
  INVX1 U13110 ( .A(n12009), .Y(n9679) );
  INVX1 U13111 ( .A(n11920), .Y(n9577) );
  INVX1 U13112 ( .A(VbeatDelay_new_1_reg_326[9]), .Y(n10474) );
  INVX1 U13113 ( .A(n11110), .Y(n10456) );
  INVX1 U13114 ( .A(ap_CS_fsm[10]), .Y(n10534) );
  AND2X1 U13115 ( .A(p_tmp_i_reg_1556[2]), .B(n8843), .Y(n8664) );
  AND2X1 U13116 ( .A(\tmp_12_reg_1694[0] ), .B(
        CircularBuffer_int_30_sum_i1_fu_1071_p3[0]), .Y(n8665) );
  AND2X1 U13117 ( .A(\tmp_s_reg_1578[0] ), .B(
        CircularBuffer_int_30_sum_i_fu_758_p3[0]), .Y(n8666) );
  INVX1 U13118 ( .A(CircularBuffer_len_read_assign_3_reg_1711[7]), .Y(n10580)
         );
  INVX1 U13119 ( .A(CircularBuffer_len_read_assign_1_reg_1616[7]), .Y(n10085)
         );
  INVX1 U13120 ( .A(recentdatapoints_head_i[0]), .Y(n9886) );
  INVX1 U13121 ( .A(n11812), .Y(n10392) );
  INVX1 U13122 ( .A(n11088), .Y(n10476) );
  INVX1 U13123 ( .A(VCaptureThresh_loc_reg_298[16]), .Y(n9705) );
  INVX1 U13124 ( .A(VCaptureThresh_loc_reg_298[20]), .Y(n9721) );
  INVX1 U13125 ( .A(ACaptureThresh_loc_reg_288[20]), .Y(n9610) );
  INVX1 U13126 ( .A(ACaptureThresh_loc_reg_288[16]), .Y(n9596) );
  INVX1 U13127 ( .A(s_axi_AXILiteS_WDATA[31]), .Y(n9282) );
  INVX1 U13128 ( .A(s_axi_AXILiteS_WDATA[30]), .Y(n9283) );
  INVX1 U13129 ( .A(s_axi_AXILiteS_WDATA[29]), .Y(n9284) );
  INVX1 U13130 ( .A(s_axi_AXILiteS_WDATA[28]), .Y(n9285) );
  INVX1 U13131 ( .A(s_axi_AXILiteS_WDATA[27]), .Y(n9286) );
  INVX1 U13132 ( .A(s_axi_AXILiteS_WDATA[26]), .Y(n9287) );
  INVX1 U13133 ( .A(s_axi_AXILiteS_WDATA[25]), .Y(n9288) );
  INVX1 U13134 ( .A(s_axi_AXILiteS_WDATA[24]), .Y(n9289) );
  INVX1 U13135 ( .A(s_axi_AXILiteS_WDATA[23]), .Y(n9290) );
  INVX1 U13136 ( .A(s_axi_AXILiteS_WDATA[22]), .Y(n9291) );
  INVX1 U13137 ( .A(s_axi_AXILiteS_WDATA[21]), .Y(n9292) );
  INVX1 U13138 ( .A(s_axi_AXILiteS_WDATA[20]), .Y(n9293) );
  INVX1 U13139 ( .A(s_axi_AXILiteS_WDATA[19]), .Y(n9294) );
  INVX1 U13140 ( .A(s_axi_AXILiteS_WDATA[18]), .Y(n9295) );
  INVX1 U13141 ( .A(s_axi_AXILiteS_WDATA[17]), .Y(n9296) );
  INVX1 U13142 ( .A(s_axi_AXILiteS_WDATA[16]), .Y(n9297) );
  INVX1 U13143 ( .A(ACaptureThresh_loc_reg_288[1]), .Y(n9550) );
  INVX1 U13144 ( .A(VCaptureThresh_loc_reg_298[1]), .Y(n9650) );
  INVX1 U13145 ( .A(CircularBuffer_len_read_assign_3_reg_1711[21]), .Y(n10594)
         );
  INVX1 U13146 ( .A(CircularBuffer_len_read_assign_1_reg_1616[21]), .Y(n10099)
         );
  AND2X1 U13147 ( .A(s_axi_AXILiteS_WVALID), .B(s_axi_AXILiteS_WREADY), .Y(
        \Decision_AXILiteS_s_axi_U/n625 ) );
  INVX1 U13148 ( .A(VbeatDelay_new_1_reg_326[13]), .Y(n10485) );
  INVX1 U13149 ( .A(VbeatDelay_new_1_reg_326[29]), .Y(n10527) );
  INVX1 U13150 ( .A(VbeatDelay_new_1_reg_326[25]), .Y(n10517) );
  INVX1 U13151 ( .A(n12051), .Y(n9719) );
  OR2X1 U13152 ( .A(n9721), .B(tmp_7_reg_1544[20]), .Y(n12050) );
  INVX1 U13153 ( .A(n12086), .Y(n9726) );
  INVX1 U13154 ( .A(n11962), .Y(n9609) );
  OR2X1 U13155 ( .A(n9610), .B(tmp_6_reg_1538[20]), .Y(n11961) );
  INVX1 U13156 ( .A(n11997), .Y(n9616) );
  INVX1 U13157 ( .A(n11854), .Y(n10419) );
  OR2X1 U13158 ( .A(n10420), .B(VbeatDelay_new_1_reg_326[20]), .Y(n11853) );
  INVX1 U13159 ( .A(n11889), .Y(n10424) );
  INVX1 U13160 ( .A(n11130), .Y(n10503) );
  OR2X1 U13161 ( .A(n10719), .B(VbeatDelay_new_1_reg_326[20]), .Y(n11129) );
  INVX1 U13162 ( .A(n11165), .Y(n10508) );
  INVX1 U13163 ( .A(CircularBuffer_len_read_assign_3_reg_1711[20]), .Y(n10593)
         );
  INVX1 U13164 ( .A(CircularBuffer_len_read_assign_3_reg_1711[6]), .Y(n10579)
         );
  INVX1 U13165 ( .A(CircularBuffer_len_read_assign_1_reg_1616[20]), .Y(n10098)
         );
  INVX1 U13166 ( .A(CircularBuffer_len_read_assign_1_reg_1616[6]), .Y(n10084)
         );
  INVX1 U13167 ( .A(AbeatDelay_new_reg_394[0]), .Y(n10677) );
  OR2X1 U13168 ( .A(n9693), .B(tmp_7_reg_1544[13]), .Y(n12018) );
  OR2X1 U13169 ( .A(n9755), .B(tmp_7_reg_1544[29]), .Y(n12065) );
  OR2X1 U13170 ( .A(n9586), .B(tmp_6_reg_1538[13]), .Y(n11929) );
  OR2X1 U13171 ( .A(n9638), .B(tmp_6_reg_1538[29]), .Y(n11976) );
  INVX1 U13172 ( .A(CircularBuffer_len_read_assign_3_reg_1711[18]), .Y(n10591)
         );
  INVX1 U13173 ( .A(CircularBuffer_len_read_assign_3_reg_1711[16]), .Y(n10589)
         );
  INVX1 U13174 ( .A(CircularBuffer_len_read_assign_3_reg_1711[12]), .Y(n10585)
         );
  INVX1 U13175 ( .A(CircularBuffer_len_read_assign_3_reg_1711[30]), .Y(n10603)
         );
  INVX1 U13176 ( .A(CircularBuffer_len_read_assign_3_reg_1711[27]), .Y(n10600)
         );
  INVX1 U13177 ( .A(CircularBuffer_len_read_assign_1_reg_1616[18]), .Y(n10096)
         );
  INVX1 U13178 ( .A(CircularBuffer_len_read_assign_1_reg_1616[16]), .Y(n10094)
         );
  INVX1 U13179 ( .A(CircularBuffer_len_read_assign_1_reg_1616[12]), .Y(n10090)
         );
  INVX1 U13180 ( .A(CircularBuffer_len_read_assign_1_reg_1616[30]), .Y(n10108)
         );
  INVX1 U13181 ( .A(CircularBuffer_len_read_assign_1_reg_1616[27]), .Y(n10105)
         );
  INVX1 U13182 ( .A(CircularBuffer_len_read_assign_3_reg_1711[17]), .Y(n10590)
         );
  INVX1 U13183 ( .A(CircularBuffer_len_read_assign_3_reg_1711[19]), .Y(n10592)
         );
  INVX1 U13184 ( .A(CircularBuffer_len_read_assign_3_reg_1711[15]), .Y(n10588)
         );
  INVX1 U13185 ( .A(CircularBuffer_len_read_assign_3_reg_1711[11]), .Y(n10584)
         );
  INVX1 U13186 ( .A(CircularBuffer_len_read_assign_3_reg_1711[26]), .Y(n10599)
         );
  INVX1 U13187 ( .A(CircularBuffer_len_read_assign_1_reg_1616[17]), .Y(n10095)
         );
  INVX1 U13188 ( .A(CircularBuffer_len_read_assign_1_reg_1616[19]), .Y(n10097)
         );
  INVX1 U13189 ( .A(CircularBuffer_len_read_assign_1_reg_1616[15]), .Y(n10093)
         );
  INVX1 U13190 ( .A(CircularBuffer_len_read_assign_1_reg_1616[11]), .Y(n10089)
         );
  INVX1 U13191 ( .A(CircularBuffer_len_read_assign_1_reg_1616[26]), .Y(n10104)
         );
  INVX1 U13192 ( .A(ap_CS_fsm[9]), .Y(n9020) );
  INVX1 U13193 ( .A(n1401), .Y(n9471) );
  INVX1 U13194 ( .A(n1515), .Y(n9496) );
  INVX1 U13195 ( .A(\Decision_AXILiteS_s_axi_U/n258 ), .Y(n9306) );
  INVX1 U13196 ( .A(\Decision_AXILiteS_s_axi_U/n265 ), .Y(n9307) );
  INVX1 U13197 ( .A(\Decision_AXILiteS_s_axi_U/n272 ), .Y(n9308) );
  INVX1 U13198 ( .A(VbeatFallDelay_new_1_reg_342[18]), .Y(n10415) );
  OR2X1 U13199 ( .A(n10401), .B(VbeatDelay_new_1_reg_326[13]), .Y(n11821) );
  OR2X1 U13200 ( .A(n10443), .B(VbeatDelay_new_1_reg_326[29]), .Y(n11868) );
  OR2X1 U13201 ( .A(n10705), .B(VbeatDelay_new_1_reg_326[13]), .Y(n11097) );
  OR2X1 U13202 ( .A(n10737), .B(VbeatDelay_new_1_reg_326[29]), .Y(n11144) );
  INVX1 U13203 ( .A(\Decision_AXILiteS_s_axi_U/n605 ), .Y(n9281) );
  OR2X1 U13204 ( .A(n10411), .B(VbeatDelay_new_1_reg_326[17]), .Y(n11879) );
  OR2X1 U13205 ( .A(n10713), .B(VbeatDelay_new_1_reg_326[17]), .Y(n11155) );
  INVX1 U13206 ( .A(n2153), .Y(n9465) );
  INVX1 U13207 ( .A(n2152), .Y(n9464) );
  INVX1 U13208 ( .A(n2151), .Y(n9463) );
  INVX1 U13209 ( .A(n2150), .Y(n9462) );
  INVX1 U13210 ( .A(n2149), .Y(n9461) );
  INVX1 U13211 ( .A(n2148), .Y(n9460) );
  INVX1 U13212 ( .A(n2147), .Y(n9459) );
  INVX1 U13213 ( .A(n2146), .Y(n9458) );
  INVX1 U13214 ( .A(n2145), .Y(n9457) );
  INVX1 U13215 ( .A(n2144), .Y(n9456) );
  INVX1 U13216 ( .A(n2143), .Y(n9455) );
  INVX1 U13217 ( .A(n2142), .Y(n9454) );
  INVX1 U13218 ( .A(n2141), .Y(n9453) );
  INVX1 U13219 ( .A(n2140), .Y(n9452) );
  INVX1 U13220 ( .A(n2139), .Y(n9451) );
  INVX1 U13221 ( .A(n2138), .Y(n9450) );
  INVX1 U13222 ( .A(n2137), .Y(n9449) );
  INVX1 U13223 ( .A(n2136), .Y(n9448) );
  INVX1 U13224 ( .A(n2135), .Y(n9447) );
  INVX1 U13225 ( .A(n2134), .Y(n9446) );
  INVX1 U13226 ( .A(n2133), .Y(n9445) );
  INVX1 U13227 ( .A(n2132), .Y(n9444) );
  INVX1 U13228 ( .A(n2131), .Y(n9443) );
  INVX1 U13229 ( .A(n2130), .Y(n9442) );
  INVX1 U13230 ( .A(n2123), .Y(n9435) );
  INVX1 U13231 ( .A(n2121), .Y(n9433) );
  INVX1 U13232 ( .A(n2120), .Y(n9432) );
  INVX1 U13233 ( .A(n2119), .Y(n9431) );
  INVX1 U13234 ( .A(n2118), .Y(n9430) );
  INVX1 U13235 ( .A(n2117), .Y(n9429) );
  INVX1 U13236 ( .A(n2116), .Y(n9428) );
  INVX1 U13237 ( .A(n2115), .Y(n9427) );
  INVX1 U13238 ( .A(n2114), .Y(n9426) );
  INVX1 U13239 ( .A(n2113), .Y(n9425) );
  INVX1 U13240 ( .A(n2112), .Y(n9424) );
  INVX1 U13241 ( .A(n2111), .Y(n9423) );
  INVX1 U13242 ( .A(n2110), .Y(n9422) );
  INVX1 U13243 ( .A(n2109), .Y(n9421) );
  INVX1 U13244 ( .A(n2108), .Y(n9420) );
  INVX1 U13245 ( .A(n2107), .Y(n9419) );
  INVX1 U13246 ( .A(n2106), .Y(n9418) );
  INVX1 U13247 ( .A(n2105), .Y(n9417) );
  INVX1 U13248 ( .A(n2104), .Y(n9416) );
  INVX1 U13249 ( .A(n2103), .Y(n9415) );
  INVX1 U13250 ( .A(n2102), .Y(n9414) );
  INVX1 U13251 ( .A(n2101), .Y(n9413) );
  INVX1 U13252 ( .A(n2100), .Y(n9412) );
  INVX1 U13253 ( .A(n2099), .Y(n9411) );
  INVX1 U13254 ( .A(n2098), .Y(n9410) );
  INVX1 U13255 ( .A(n2097), .Y(n9409) );
  INVX1 U13256 ( .A(n2093), .Y(n9405) );
  INVX1 U13257 ( .A(n2092), .Y(n9404) );
  INVX1 U13258 ( .A(n2129), .Y(n9441) );
  INVX1 U13259 ( .A(n2128), .Y(n9440) );
  INVX1 U13260 ( .A(n2127), .Y(n9439) );
  INVX1 U13261 ( .A(n2126), .Y(n9438) );
  INVX1 U13262 ( .A(n2125), .Y(n9437) );
  INVX1 U13263 ( .A(n2124), .Y(n9436) );
  INVX1 U13264 ( .A(n2122), .Y(n9434) );
  INVX1 U13265 ( .A(n2096), .Y(n9408) );
  INVX1 U13266 ( .A(n2095), .Y(n9407) );
  INVX1 U13267 ( .A(n2094), .Y(n9406) );
  INVX1 U13268 ( .A(n2091), .Y(n9403) );
  INVX1 U13269 ( .A(n2088), .Y(n9402) );
  INVX1 U13270 ( .A(VbeatFallDelay_new_1_reg_342[24]), .Y(n10431) );
  INVX1 U13271 ( .A(VbeatFallDelay_new_1_reg_342[2]), .Y(n10373) );
  INVX1 U13272 ( .A(VbeatFallDelay_new_1_reg_342[26]), .Y(n10437) );
  INVX1 U13273 ( .A(VbeatFallDelay_new_1_reg_342[30]), .Y(n10447) );
  OR2X1 U13274 ( .A(n9741), .B(tmp_7_reg_1544[25]), .Y(n12058) );
  OR2X1 U13275 ( .A(n9626), .B(tmp_6_reg_1538[25]), .Y(n11969) );
  INVX1 U13276 ( .A(VbeatFallDelay_new_1_reg_342[6]), .Y(n10382) );
  INVX1 U13277 ( .A(VbeatFallDelay_new_1_reg_342[14]), .Y(n10405) );
  INVX1 U13278 ( .A(VbeatFallDelay_new_1_reg_342[22]), .Y(n10426) );
  INVX1 U13279 ( .A(VbeatFallDelay_new_1_reg_342[17]), .Y(n10411) );
  INVX1 U13280 ( .A(n2071), .Y(n9386) );
  INVX1 U13281 ( .A(n2073), .Y(n9387) );
  INVX1 U13282 ( .A(n2074), .Y(n9388) );
  INVX1 U13283 ( .A(n2075), .Y(n9389) );
  INVX1 U13284 ( .A(n2076), .Y(n9390) );
  INVX1 U13285 ( .A(n2077), .Y(n9391) );
  INVX1 U13286 ( .A(n2078), .Y(n9392) );
  INVX1 U13287 ( .A(n2079), .Y(n9393) );
  INVX1 U13288 ( .A(n2080), .Y(n9394) );
  INVX1 U13289 ( .A(n2081), .Y(n9395) );
  INVX1 U13290 ( .A(n2082), .Y(n9396) );
  INVX1 U13291 ( .A(n2083), .Y(n9397) );
  INVX1 U13292 ( .A(n2084), .Y(n9398) );
  INVX1 U13293 ( .A(n2085), .Y(n9399) );
  INVX1 U13294 ( .A(n2086), .Y(n9400) );
  INVX1 U13295 ( .A(n2087), .Y(n9401) );
  OR2X1 U13296 ( .A(n9707), .B(tmp_7_reg_1544[17]), .Y(n12076) );
  OR2X1 U13297 ( .A(n9724), .B(tmp_7_reg_1544[21]), .Y(n12083) );
  OR2X1 U13298 ( .A(n9598), .B(tmp_6_reg_1538[17]), .Y(n11987) );
  OR2X1 U13299 ( .A(n9612), .B(tmp_6_reg_1538[21]), .Y(n11994) );
  INVX1 U13300 ( .A(recentABools_sum[0]), .Y(n10543) );
  INVX1 U13301 ( .A(recentVBools_sum[0]), .Y(n10208) );
  INVX1 U13302 ( .A(recentABools_sum[1]), .Y(n10544) );
  INVX1 U13303 ( .A(recentVBools_sum[1]), .Y(n10209) );
  INVX1 U13304 ( .A(recentABools_sum[2]), .Y(n10545) );
  INVX1 U13305 ( .A(recentVBools_sum[2]), .Y(n10210) );
  INVX1 U13306 ( .A(recentABools_sum[3]), .Y(n10546) );
  INVX1 U13307 ( .A(recentVBools_sum[3]), .Y(n10211) );
  INVX1 U13308 ( .A(recentABools_sum[4]), .Y(n10547) );
  INVX1 U13309 ( .A(recentVBools_sum[4]), .Y(n10212) );
  INVX1 U13310 ( .A(recentABools_sum[5]), .Y(n10548) );
  INVX1 U13311 ( .A(recentVBools_sum[5]), .Y(n10213) );
  INVX1 U13312 ( .A(recentABools_sum[6]), .Y(n10549) );
  INVX1 U13313 ( .A(recentVBools_sum[6]), .Y(n10214) );
  INVX1 U13314 ( .A(recentABools_sum[7]), .Y(n10550) );
  INVX1 U13315 ( .A(recentVBools_sum[7]), .Y(n10215) );
  INVX1 U13316 ( .A(recentABools_sum[8]), .Y(n10551) );
  INVX1 U13317 ( .A(recentVBools_sum[8]), .Y(n10216) );
  INVX1 U13318 ( .A(recentABools_sum[9]), .Y(n10552) );
  INVX1 U13319 ( .A(recentVBools_sum[9]), .Y(n10217) );
  INVX1 U13320 ( .A(recentABools_sum[10]), .Y(n10553) );
  INVX1 U13321 ( .A(recentVBools_sum[10]), .Y(n10218) );
  INVX1 U13322 ( .A(recentABools_sum[11]), .Y(n10554) );
  INVX1 U13323 ( .A(recentVBools_sum[11]), .Y(n10219) );
  INVX1 U13324 ( .A(recentABools_sum[12]), .Y(n10555) );
  INVX1 U13325 ( .A(recentVBools_sum[12]), .Y(n10220) );
  INVX1 U13326 ( .A(recentABools_sum[13]), .Y(n10556) );
  INVX1 U13327 ( .A(recentVBools_sum[13]), .Y(n10221) );
  INVX1 U13328 ( .A(recentABools_sum[14]), .Y(n10557) );
  INVX1 U13329 ( .A(recentVBools_sum[14]), .Y(n10222) );
  INVX1 U13330 ( .A(recentABools_sum[15]), .Y(n10558) );
  INVX1 U13331 ( .A(recentVBools_sum[15]), .Y(n10223) );
  INVX1 U13332 ( .A(recentABools_sum[16]), .Y(n10559) );
  INVX1 U13333 ( .A(recentVBools_sum[16]), .Y(n10224) );
  INVX1 U13334 ( .A(recentABools_sum[17]), .Y(n10560) );
  INVX1 U13335 ( .A(recentVBools_sum[17]), .Y(n10225) );
  INVX1 U13336 ( .A(recentABools_sum[18]), .Y(n10561) );
  INVX1 U13337 ( .A(recentVBools_sum[18]), .Y(n10226) );
  INVX1 U13338 ( .A(recentABools_sum[19]), .Y(n10562) );
  INVX1 U13339 ( .A(recentVBools_sum[19]), .Y(n10227) );
  INVX1 U13340 ( .A(recentABools_sum[20]), .Y(n10563) );
  INVX1 U13341 ( .A(recentVBools_sum[20]), .Y(n10228) );
  INVX1 U13342 ( .A(recentABools_sum[21]), .Y(n10564) );
  INVX1 U13343 ( .A(recentVBools_sum[21]), .Y(n10229) );
  INVX1 U13344 ( .A(recentABools_sum[22]), .Y(n10565) );
  INVX1 U13345 ( .A(recentVBools_sum[22]), .Y(n10230) );
  INVX1 U13346 ( .A(recentABools_sum[23]), .Y(n10566) );
  INVX1 U13347 ( .A(recentVBools_sum[23]), .Y(n10231) );
  INVX1 U13348 ( .A(recentABools_sum[24]), .Y(n10567) );
  INVX1 U13349 ( .A(recentVBools_sum[24]), .Y(n10232) );
  INVX1 U13350 ( .A(recentABools_sum[25]), .Y(n10568) );
  INVX1 U13351 ( .A(recentVBools_sum[25]), .Y(n10233) );
  INVX1 U13352 ( .A(recentABools_sum[26]), .Y(n10569) );
  INVX1 U13353 ( .A(recentVBools_sum[26]), .Y(n10234) );
  INVX1 U13354 ( .A(recentABools_sum[27]), .Y(n10570) );
  INVX1 U13355 ( .A(recentVBools_sum[27]), .Y(n10235) );
  INVX1 U13356 ( .A(recentABools_sum[28]), .Y(n10571) );
  INVX1 U13357 ( .A(recentVBools_sum[28]), .Y(n10236) );
  INVX1 U13358 ( .A(recentABools_sum[29]), .Y(n10572) );
  INVX1 U13359 ( .A(recentVBools_sum[29]), .Y(n10237) );
  INVX1 U13360 ( .A(recentABools_sum[30]), .Y(n10811) );
  INVX1 U13361 ( .A(recentVBools_sum[30]), .Y(n10238) );
  INVX1 U13362 ( .A(VbeatFallDelay_new_1_reg_342[12]), .Y(n10399) );
  INVX1 U13363 ( .A(VbeatFallDelay_new_1_reg_342[28]), .Y(n10441) );
  INVX1 U13364 ( .A(VbeatDelay_new_1_reg_326[0]), .Y(n10451) );
  INVX1 U13365 ( .A(VbeatFallDelay_new_1_reg_342[5]), .Y(n10379) );
  INVX1 U13366 ( .A(VbeatFallDelay_new_1_reg_342[1]), .Y(n10370) );
  OR2X1 U13367 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[0]), .B(n10667), 
        .Y(n8667) );
  OR2X1 U13368 ( .A(CircularBuffer_sum_read_assign_reg_1610[0]), .B(n10207), 
        .Y(n8668) );
  OR2X1 U13369 ( .A(recentABools_sum[0]), .B(n10666), .Y(n8669) );
  OR2X1 U13370 ( .A(recentVBools_sum[0]), .B(n10206), .Y(n8670) );
  OR2X1 U13371 ( .A(n10422), .B(VbeatDelay_new_1_reg_326[21]), .Y(n11886) );
  OR2X1 U13372 ( .A(n10721), .B(VbeatDelay_new_1_reg_326[21]), .Y(n11162) );
  OR2X1 U13373 ( .A(n10433), .B(VbeatDelay_new_1_reg_326[25]), .Y(n11861) );
  OR2X1 U13374 ( .A(n10729), .B(VbeatDelay_new_1_reg_326[25]), .Y(n11137) );
  OR2X1 U13375 ( .A(CircularBuffer_len_read_assign_3_reg_1711[3]), .B(n8841), 
        .Y(n8671) );
  OR2X1 U13376 ( .A(CircularBuffer_len_read_assign_1_reg_1616[3]), .B(n8842), 
        .Y(n8672) );
  INVX1 U13377 ( .A(CircularBuffer_len_write_assig_2_reg_1729[5]), .Y(n10639)
         );
  INVX1 U13378 ( .A(CircularBuffer_len_write_assig_reg_1634[5]), .Y(n10144) );
  OR2X1 U13379 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[2]), .B(n8837), 
        .Y(n8673) );
  OR2X1 U13380 ( .A(CircularBuffer_sum_read_assign_reg_1610[2]), .B(n8838), 
        .Y(n8674) );
  OR2X1 U13381 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[3]), .B(n8673), 
        .Y(n8675) );
  OR2X1 U13382 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[4]), .B(n8675), 
        .Y(n8676) );
  OR2X1 U13383 ( .A(CircularBuffer_sum_read_assign_reg_1610[3]), .B(n8674), 
        .Y(n8677) );
  OR2X1 U13384 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[5]), .B(n8676), 
        .Y(n8678) );
  OR2X1 U13385 ( .A(CircularBuffer_sum_read_assign_reg_1610[4]), .B(n8677), 
        .Y(n8679) );
  OR2X1 U13386 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[6]), .B(n8678), 
        .Y(n8680) );
  OR2X1 U13387 ( .A(CircularBuffer_sum_read_assign_reg_1610[5]), .B(n8679), 
        .Y(n8681) );
  OR2X1 U13388 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[7]), .B(n8680), 
        .Y(n8682) );
  OR2X1 U13389 ( .A(CircularBuffer_sum_read_assign_reg_1610[6]), .B(n8681), 
        .Y(n8683) );
  OR2X1 U13390 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[8]), .B(n8682), 
        .Y(n8684) );
  OR2X1 U13391 ( .A(CircularBuffer_sum_read_assign_reg_1610[7]), .B(n8683), 
        .Y(n8685) );
  OR2X1 U13392 ( .A(recentABools_sum[2]), .B(n8839), .Y(n8686) );
  OR2X1 U13393 ( .A(recentVBools_sum[2]), .B(n8840), .Y(n8687) );
  OR2X1 U13394 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[9]), .B(n8684), 
        .Y(n8688) );
  OR2X1 U13395 ( .A(CircularBuffer_sum_read_assign_reg_1610[8]), .B(n8685), 
        .Y(n8689) );
  OR2X1 U13396 ( .A(recentABools_sum[3]), .B(n8686), .Y(n8690) );
  OR2X1 U13397 ( .A(recentVBools_sum[3]), .B(n8687), .Y(n8691) );
  OR2X1 U13398 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[10]), .B(n8688), 
        .Y(n8692) );
  OR2X1 U13399 ( .A(CircularBuffer_sum_read_assign_reg_1610[9]), .B(n8689), 
        .Y(n8693) );
  OR2X1 U13400 ( .A(recentABools_sum[4]), .B(n8690), .Y(n8694) );
  OR2X1 U13401 ( .A(recentVBools_sum[4]), .B(n8691), .Y(n8695) );
  OR2X1 U13402 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[11]), .B(n8692), 
        .Y(n8696) );
  OR2X1 U13403 ( .A(CircularBuffer_sum_read_assign_reg_1610[10]), .B(n8693), 
        .Y(n8697) );
  OR2X1 U13404 ( .A(recentABools_sum[5]), .B(n8694), .Y(n8698) );
  OR2X1 U13405 ( .A(recentVBools_sum[5]), .B(n8695), .Y(n8699) );
  OR2X1 U13406 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[12]), .B(n8696), 
        .Y(n8700) );
  OR2X1 U13407 ( .A(CircularBuffer_sum_read_assign_reg_1610[11]), .B(n8697), 
        .Y(n8701) );
  OR2X1 U13408 ( .A(recentABools_sum[6]), .B(n8698), .Y(n8702) );
  OR2X1 U13409 ( .A(recentVBools_sum[6]), .B(n8699), .Y(n8703) );
  OR2X1 U13410 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[13]), .B(n8700), 
        .Y(n8704) );
  OR2X1 U13411 ( .A(CircularBuffer_len_read_assign_3_reg_1711[5]), .B(n8835), 
        .Y(n8705) );
  OR2X1 U13412 ( .A(CircularBuffer_sum_read_assign_reg_1610[12]), .B(n8701), 
        .Y(n8706) );
  OR2X1 U13413 ( .A(CircularBuffer_len_read_assign_1_reg_1616[5]), .B(n8836), 
        .Y(n8707) );
  OR2X1 U13414 ( .A(recentABools_sum[7]), .B(n8702), .Y(n8708) );
  OR2X1 U13415 ( .A(recentVBools_sum[7]), .B(n8703), .Y(n8709) );
  OR2X1 U13416 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[14]), .B(n8704), 
        .Y(n8710) );
  OR2X1 U13417 ( .A(CircularBuffer_len_read_assign_3_reg_1711[6]), .B(n8705), 
        .Y(n8711) );
  OR2X1 U13418 ( .A(CircularBuffer_sum_read_assign_reg_1610[13]), .B(n8706), 
        .Y(n8712) );
  OR2X1 U13419 ( .A(CircularBuffer_len_read_assign_1_reg_1616[6]), .B(n8707), 
        .Y(n8713) );
  OR2X1 U13420 ( .A(recentABools_sum[8]), .B(n8708), .Y(n8714) );
  OR2X1 U13421 ( .A(recentVBools_sum[8]), .B(n8709), .Y(n8715) );
  OR2X1 U13422 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[15]), .B(n8710), 
        .Y(n8716) );
  OR2X1 U13423 ( .A(CircularBuffer_len_read_assign_3_reg_1711[7]), .B(n8711), 
        .Y(n8717) );
  OR2X1 U13424 ( .A(CircularBuffer_sum_read_assign_reg_1610[14]), .B(n8712), 
        .Y(n8718) );
  OR2X1 U13425 ( .A(CircularBuffer_len_read_assign_1_reg_1616[7]), .B(n8713), 
        .Y(n8719) );
  OR2X1 U13426 ( .A(recentABools_sum[9]), .B(n8714), .Y(n8720) );
  OR2X1 U13427 ( .A(recentVBools_sum[9]), .B(n8715), .Y(n8721) );
  OR2X1 U13428 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[16]), .B(n8716), 
        .Y(n8722) );
  OR2X1 U13429 ( .A(CircularBuffer_len_read_assign_3_reg_1711[8]), .B(n8717), 
        .Y(n8723) );
  OR2X1 U13430 ( .A(CircularBuffer_sum_read_assign_reg_1610[15]), .B(n8718), 
        .Y(n8724) );
  OR2X1 U13431 ( .A(CircularBuffer_len_read_assign_1_reg_1616[8]), .B(n8719), 
        .Y(n8725) );
  OR2X1 U13432 ( .A(recentABools_sum[10]), .B(n8720), .Y(n8726) );
  OR2X1 U13433 ( .A(recentVBools_sum[10]), .B(n8721), .Y(n8727) );
  OR2X1 U13434 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[17]), .B(n8722), 
        .Y(n8728) );
  OR2X1 U13435 ( .A(CircularBuffer_len_read_assign_3_reg_1711[9]), .B(n8723), 
        .Y(n8729) );
  OR2X1 U13436 ( .A(CircularBuffer_sum_read_assign_reg_1610[16]), .B(n8724), 
        .Y(n8730) );
  OR2X1 U13437 ( .A(CircularBuffer_len_read_assign_1_reg_1616[9]), .B(n8725), 
        .Y(n8731) );
  OR2X1 U13438 ( .A(recentABools_sum[11]), .B(n8726), .Y(n8732) );
  OR2X1 U13439 ( .A(recentVBools_sum[11]), .B(n8727), .Y(n8733) );
  OR2X1 U13440 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[18]), .B(n8728), 
        .Y(n8734) );
  OR2X1 U13441 ( .A(CircularBuffer_len_read_assign_3_reg_1711[10]), .B(n8729), 
        .Y(n8735) );
  OR2X1 U13442 ( .A(CircularBuffer_sum_read_assign_reg_1610[17]), .B(n8730), 
        .Y(n8736) );
  OR2X1 U13443 ( .A(CircularBuffer_len_read_assign_1_reg_1616[10]), .B(n8731), 
        .Y(n8737) );
  OR2X1 U13444 ( .A(recentABools_sum[12]), .B(n8732), .Y(n8738) );
  OR2X1 U13445 ( .A(recentVBools_sum[12]), .B(n8733), .Y(n8739) );
  OR2X1 U13446 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[19]), .B(n8734), 
        .Y(n8740) );
  OR2X1 U13447 ( .A(CircularBuffer_len_read_assign_3_reg_1711[11]), .B(n8735), 
        .Y(n8741) );
  OR2X1 U13448 ( .A(CircularBuffer_sum_read_assign_reg_1610[18]), .B(n8736), 
        .Y(n8742) );
  OR2X1 U13449 ( .A(CircularBuffer_len_read_assign_1_reg_1616[11]), .B(n8737), 
        .Y(n8743) );
  OR2X1 U13450 ( .A(recentABools_sum[13]), .B(n8738), .Y(n8744) );
  OR2X1 U13451 ( .A(recentVBools_sum[13]), .B(n8739), .Y(n8745) );
  OR2X1 U13452 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[20]), .B(n8740), 
        .Y(n8746) );
  OR2X1 U13453 ( .A(CircularBuffer_len_read_assign_3_reg_1711[12]), .B(n8741), 
        .Y(n8747) );
  OR2X1 U13454 ( .A(CircularBuffer_sum_read_assign_reg_1610[19]), .B(n8742), 
        .Y(n8748) );
  OR2X1 U13455 ( .A(CircularBuffer_len_read_assign_1_reg_1616[12]), .B(n8743), 
        .Y(n8749) );
  OR2X1 U13456 ( .A(recentABools_sum[14]), .B(n8744), .Y(n8750) );
  OR2X1 U13457 ( .A(recentVBools_sum[14]), .B(n8745), .Y(n8751) );
  OR2X1 U13458 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[21]), .B(n8746), 
        .Y(n8752) );
  OR2X1 U13459 ( .A(CircularBuffer_len_read_assign_3_reg_1711[13]), .B(n8747), 
        .Y(n8753) );
  OR2X1 U13460 ( .A(CircularBuffer_sum_read_assign_reg_1610[20]), .B(n8748), 
        .Y(n8754) );
  OR2X1 U13461 ( .A(CircularBuffer_len_read_assign_1_reg_1616[13]), .B(n8749), 
        .Y(n8755) );
  OR2X1 U13462 ( .A(recentABools_sum[15]), .B(n8750), .Y(n8756) );
  OR2X1 U13463 ( .A(recentVBools_sum[15]), .B(n8751), .Y(n8757) );
  OR2X1 U13464 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[22]), .B(n8752), 
        .Y(n8758) );
  OR2X1 U13465 ( .A(CircularBuffer_len_read_assign_3_reg_1711[14]), .B(n8753), 
        .Y(n8759) );
  OR2X1 U13466 ( .A(CircularBuffer_sum_read_assign_reg_1610[21]), .B(n8754), 
        .Y(n8760) );
  OR2X1 U13467 ( .A(CircularBuffer_len_read_assign_1_reg_1616[14]), .B(n8755), 
        .Y(n8761) );
  OR2X1 U13468 ( .A(recentABools_sum[16]), .B(n8756), .Y(n8762) );
  OR2X1 U13469 ( .A(recentVBools_sum[16]), .B(n8757), .Y(n8763) );
  OR2X1 U13470 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[23]), .B(n8758), 
        .Y(n8764) );
  OR2X1 U13471 ( .A(CircularBuffer_len_read_assign_3_reg_1711[15]), .B(n8759), 
        .Y(n8765) );
  OR2X1 U13472 ( .A(CircularBuffer_sum_read_assign_reg_1610[22]), .B(n8760), 
        .Y(n8766) );
  OR2X1 U13473 ( .A(CircularBuffer_len_read_assign_1_reg_1616[15]), .B(n8761), 
        .Y(n8767) );
  OR2X1 U13474 ( .A(recentABools_sum[17]), .B(n8762), .Y(n8768) );
  OR2X1 U13475 ( .A(recentVBools_sum[17]), .B(n8763), .Y(n8769) );
  OR2X1 U13476 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[24]), .B(n8764), 
        .Y(n8770) );
  OR2X1 U13477 ( .A(CircularBuffer_len_read_assign_3_reg_1711[16]), .B(n8765), 
        .Y(n8771) );
  OR2X1 U13478 ( .A(CircularBuffer_sum_read_assign_reg_1610[23]), .B(n8766), 
        .Y(n8772) );
  OR2X1 U13479 ( .A(CircularBuffer_len_read_assign_1_reg_1616[16]), .B(n8767), 
        .Y(n8773) );
  OR2X1 U13480 ( .A(recentABools_sum[18]), .B(n8768), .Y(n8774) );
  OR2X1 U13481 ( .A(recentVBools_sum[18]), .B(n8769), .Y(n8775) );
  OR2X1 U13482 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[25]), .B(n8770), 
        .Y(n8776) );
  OR2X1 U13483 ( .A(CircularBuffer_len_read_assign_3_reg_1711[17]), .B(n8771), 
        .Y(n8777) );
  OR2X1 U13484 ( .A(CircularBuffer_sum_read_assign_reg_1610[24]), .B(n8772), 
        .Y(n8778) );
  OR2X1 U13485 ( .A(CircularBuffer_len_read_assign_1_reg_1616[17]), .B(n8773), 
        .Y(n8779) );
  OR2X1 U13486 ( .A(recentABools_sum[19]), .B(n8774), .Y(n8780) );
  OR2X1 U13487 ( .A(recentVBools_sum[19]), .B(n8775), .Y(n8781) );
  OR2X1 U13488 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[26]), .B(n8776), 
        .Y(n8782) );
  OR2X1 U13489 ( .A(CircularBuffer_len_read_assign_3_reg_1711[18]), .B(n8777), 
        .Y(n8783) );
  OR2X1 U13490 ( .A(CircularBuffer_sum_read_assign_reg_1610[25]), .B(n8778), 
        .Y(n8784) );
  OR2X1 U13491 ( .A(CircularBuffer_len_read_assign_1_reg_1616[18]), .B(n8779), 
        .Y(n8785) );
  OR2X1 U13492 ( .A(recentABools_sum[20]), .B(n8780), .Y(n8786) );
  OR2X1 U13493 ( .A(recentVBools_sum[20]), .B(n8781), .Y(n8787) );
  OR2X1 U13494 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[27]), .B(n8782), 
        .Y(n8788) );
  OR2X1 U13495 ( .A(CircularBuffer_len_read_assign_3_reg_1711[19]), .B(n8783), 
        .Y(n8789) );
  OR2X1 U13496 ( .A(CircularBuffer_sum_read_assign_reg_1610[26]), .B(n8784), 
        .Y(n8790) );
  OR2X1 U13497 ( .A(CircularBuffer_len_read_assign_1_reg_1616[19]), .B(n8785), 
        .Y(n8791) );
  OR2X1 U13498 ( .A(recentABools_sum[21]), .B(n8786), .Y(n8792) );
  OR2X1 U13499 ( .A(recentVBools_sum[21]), .B(n8787), .Y(n8793) );
  OR2X1 U13500 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[28]), .B(n8788), 
        .Y(n8794) );
  OR2X1 U13501 ( .A(CircularBuffer_len_read_assign_3_reg_1711[20]), .B(n8789), 
        .Y(n8795) );
  OR2X1 U13502 ( .A(CircularBuffer_sum_read_assign_reg_1610[27]), .B(n8790), 
        .Y(n8796) );
  OR2X1 U13503 ( .A(CircularBuffer_len_read_assign_1_reg_1616[20]), .B(n8791), 
        .Y(n8797) );
  OR2X1 U13504 ( .A(recentABools_sum[22]), .B(n8792), .Y(n8798) );
  OR2X1 U13505 ( .A(recentVBools_sum[22]), .B(n8793), .Y(n8799) );
  OR2X1 U13506 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[29]), .B(n8794), 
        .Y(n8800) );
  OR2X1 U13507 ( .A(CircularBuffer_len_read_assign_3_reg_1711[21]), .B(n8795), 
        .Y(n8801) );
  OR2X1 U13508 ( .A(CircularBuffer_sum_read_assign_reg_1610[28]), .B(n8796), 
        .Y(n8802) );
  OR2X1 U13509 ( .A(CircularBuffer_len_read_assign_1_reg_1616[21]), .B(n8797), 
        .Y(n8803) );
  OR2X1 U13510 ( .A(recentABools_sum[23]), .B(n8798), .Y(n8804) );
  OR2X1 U13511 ( .A(recentVBools_sum[23]), .B(n8799), .Y(n8805) );
  OR2X1 U13512 ( .A(CircularBuffer_len_read_assign_3_reg_1711[22]), .B(n8801), 
        .Y(n8806) );
  OR2X1 U13513 ( .A(CircularBuffer_sum_read_assign_reg_1610[29]), .B(n8802), 
        .Y(n8807) );
  OR2X1 U13514 ( .A(CircularBuffer_len_read_assign_1_reg_1616[22]), .B(n8803), 
        .Y(n8808) );
  OR2X1 U13515 ( .A(recentABools_sum[24]), .B(n8804), .Y(n8809) );
  OR2X1 U13516 ( .A(recentVBools_sum[24]), .B(n8805), .Y(n8810) );
  OR2X1 U13517 ( .A(CircularBuffer_len_read_assign_3_reg_1711[23]), .B(n8806), 
        .Y(n8811) );
  OR2X1 U13518 ( .A(CircularBuffer_len_read_assign_1_reg_1616[23]), .B(n8808), 
        .Y(n8812) );
  OR2X1 U13519 ( .A(recentABools_sum[25]), .B(n8809), .Y(n8813) );
  OR2X1 U13520 ( .A(recentVBools_sum[25]), .B(n8810), .Y(n8814) );
  OR2X1 U13521 ( .A(CircularBuffer_len_read_assign_3_reg_1711[24]), .B(n8811), 
        .Y(n8815) );
  OR2X1 U13522 ( .A(CircularBuffer_len_read_assign_1_reg_1616[24]), .B(n8812), 
        .Y(n8816) );
  OR2X1 U13523 ( .A(recentABools_sum[26]), .B(n8813), .Y(n8817) );
  OR2X1 U13524 ( .A(recentVBools_sum[26]), .B(n8814), .Y(n8818) );
  OR2X1 U13525 ( .A(CircularBuffer_len_read_assign_3_reg_1711[25]), .B(n8815), 
        .Y(n8819) );
  OR2X1 U13526 ( .A(CircularBuffer_len_read_assign_1_reg_1616[25]), .B(n8816), 
        .Y(n8820) );
  OR2X1 U13527 ( .A(recentABools_sum[27]), .B(n8817), .Y(n8821) );
  OR2X1 U13528 ( .A(recentVBools_sum[27]), .B(n8818), .Y(n8822) );
  OR2X1 U13529 ( .A(CircularBuffer_len_read_assign_3_reg_1711[26]), .B(n8819), 
        .Y(n8823) );
  OR2X1 U13530 ( .A(CircularBuffer_len_read_assign_1_reg_1616[26]), .B(n8820), 
        .Y(n8824) );
  OR2X1 U13531 ( .A(recentABools_sum[28]), .B(n8821), .Y(n8825) );
  OR2X1 U13532 ( .A(recentVBools_sum[28]), .B(n8822), .Y(n8826) );
  OR2X1 U13533 ( .A(CircularBuffer_len_read_assign_3_reg_1711[27]), .B(n8823), 
        .Y(n8827) );
  OR2X1 U13534 ( .A(CircularBuffer_len_read_assign_1_reg_1616[27]), .B(n8824), 
        .Y(n8828) );
  OR2X1 U13535 ( .A(recentABools_sum[29]), .B(n8825), .Y(n8829) );
  OR2X1 U13536 ( .A(recentVBools_sum[29]), .B(n8826), .Y(n8830) );
  OR2X1 U13537 ( .A(CircularBuffer_len_read_assign_3_reg_1711[28]), .B(n8827), 
        .Y(n8831) );
  OR2X1 U13538 ( .A(CircularBuffer_len_read_assign_1_reg_1616[28]), .B(n8828), 
        .Y(n8832) );
  OR2X1 U13539 ( .A(CircularBuffer_len_read_assign_3_reg_1711[29]), .B(n8831), 
        .Y(n8833) );
  OR2X1 U13540 ( .A(CircularBuffer_len_read_assign_1_reg_1616[29]), .B(n8832), 
        .Y(n8834) );
  OR2X1 U13541 ( .A(CircularBuffer_len_read_assign_3_reg_1711[4]), .B(n8671), 
        .Y(n8835) );
  OR2X1 U13542 ( .A(CircularBuffer_len_read_assign_1_reg_1616[4]), .B(n8672), 
        .Y(n8836) );
  OR2X1 U13543 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[1]), .B(n8667), 
        .Y(n8837) );
  OR2X1 U13544 ( .A(CircularBuffer_sum_read_assign_reg_1610[1]), .B(n8668), 
        .Y(n8838) );
  OR2X1 U13545 ( .A(recentABools_sum[1]), .B(n8669), .Y(n8839) );
  OR2X1 U13546 ( .A(recentVBools_sum[1]), .B(n8670), .Y(n8840) );
  INVX1 U13547 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[8]), .Y(n10334)
         );
  INVX1 U13548 ( .A(CircularBuffer_head_i_read_ass_reg_1624[8]), .Y(n10027) );
  INVX1 U13549 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[10]), .Y(n10336)
         );
  INVX1 U13550 ( .A(CircularBuffer_head_i_read_ass_reg_1624[10]), .Y(n10029)
         );
  INVX1 U13551 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[12]), .Y(n10338)
         );
  INVX1 U13552 ( .A(CircularBuffer_head_i_read_ass_reg_1624[12]), .Y(n10031)
         );
  INVX1 U13553 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[14]), .Y(n10340)
         );
  INVX1 U13554 ( .A(CircularBuffer_head_i_read_ass_reg_1624[14]), .Y(n10033)
         );
  INVX1 U13555 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[16]), .Y(n10342)
         );
  INVX1 U13556 ( .A(CircularBuffer_head_i_read_ass_reg_1624[16]), .Y(n10035)
         );
  INVX1 U13557 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[18]), .Y(n10344)
         );
  INVX1 U13558 ( .A(CircularBuffer_head_i_read_ass_reg_1624[18]), .Y(n10037)
         );
  INVX1 U13559 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[20]), .Y(n10346)
         );
  INVX1 U13560 ( .A(CircularBuffer_head_i_read_ass_reg_1624[20]), .Y(n10039)
         );
  INVX1 U13561 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[22]), .Y(n10348)
         );
  INVX1 U13562 ( .A(CircularBuffer_head_i_read_ass_reg_1624[22]), .Y(n10041)
         );
  INVX1 U13563 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[24]), .Y(n10350)
         );
  INVX1 U13564 ( .A(CircularBuffer_head_i_read_ass_reg_1624[24]), .Y(n10043)
         );
  INVX1 U13565 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[26]), .Y(n10352)
         );
  INVX1 U13566 ( .A(CircularBuffer_head_i_read_ass_reg_1624[26]), .Y(n10045)
         );
  INVX1 U13567 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[28]), .Y(n10354)
         );
  INVX1 U13568 ( .A(CircularBuffer_head_i_read_ass_reg_1624[28]), .Y(n10047)
         );
  INVX1 U13569 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[29]), .Y(n10355)
         );
  INVX1 U13570 ( .A(CircularBuffer_head_i_read_ass_reg_1624[29]), .Y(n10048)
         );
  INVX1 U13571 ( .A(VbeatFallDelay_new_1_reg_342[21]), .Y(n10422) );
  INVX1 U13572 ( .A(VbeatFallDelay_new_1_reg_342[4]), .Y(n10377) );
  INVX1 U13573 ( .A(ap_CS_fsm[8]), .Y(n10242) );
  INVX1 U13574 ( .A(ap_CS_fsm[3]), .Y(n9934) );
  AND2X1 U13575 ( .A(\Decision_AXILiteS_s_axi_U/wstate[0] ), .B(n10900), .Y(
        s_axi_AXILiteS_WREADY) );
  INVX1 U13576 ( .A(\Decision_AXILiteS_s_axi_U/int_isr[0] ), .Y(n10885) );
  INVX1 U13577 ( .A(tmp_7_reg_1544[1]), .Y(n10778) );
  INVX1 U13578 ( .A(tmp_6_reg_1538[1]), .Y(n10744) );
  INVX1 U13579 ( .A(VbeatFallDelay_new_1_reg_342[9]), .Y(n10390) );
  INVX1 U13580 ( .A(VbeatFallDelay_new_1_reg_342[16]), .Y(n10409) );
  OR2X1 U13581 ( .A(CircularBuffer_len_read_assign_3_reg_1711[2]), .B(
        CircularBuffer_len_read_assign_3_reg_1711[1]), .Y(n8841) );
  OR2X1 U13582 ( .A(CircularBuffer_len_read_assign_1_reg_1616[2]), .B(
        CircularBuffer_len_read_assign_1_reg_1616[1]), .Y(n8842) );
  OR2X1 U13583 ( .A(n9661), .B(tmp_7_reg_1544[5]), .Y(n12039) );
  OR2X1 U13584 ( .A(n9560), .B(tmp_6_reg_1538[5]), .Y(n11950) );
  OR2X1 U13585 ( .A(p_tmp_i_reg_1556[1]), .B(p_tmp_i_reg_1556[0]), .Y(n8843)
         );
  INVX1 U13586 ( .A(VbeatFallDelay_new_1_reg_342[13]), .Y(n10401) );
  INVX1 U13587 ( .A(VbeatFallDelay_new_1_reg_342[29]), .Y(n10443) );
  INVX1 U13588 ( .A(VbeatFallDelay_new_1_reg_342[25]), .Y(n10433) );
  INVX1 U13589 ( .A(recentABools_len[0]), .Y(n10540) );
  INVX1 U13590 ( .A(recentVBools_len[0]), .Y(n10075) );
  INVX1 U13591 ( .A(ap_CS_fsm[6]), .Y(n10057) );
  INVX1 U13592 ( .A(ap_CS_fsm[11]), .Y(n10535) );
  INVX1 U13593 ( .A(VbeatFallDelay_new_1_reg_342[20]), .Y(n10420) );
  OR2X1 U13594 ( .A(n10379), .B(VbeatDelay_new_1_reg_326[5]), .Y(n11842) );
  OR2X1 U13595 ( .A(n10689), .B(VbeatDelay_new_1_reg_326[5]), .Y(n11118) );
  INVX1 U13596 ( .A(tmp_7_reg_1544[24]), .Y(n10801) );
  INVX1 U13597 ( .A(tmp_6_reg_1538[24]), .Y(n10767) );
  INVX1 U13598 ( .A(tmp_38_i_reg_1550[7]), .Y(n9925) );
  AND2X1 U13599 ( .A(ap_CS_fsm[2]), .B(ap_rst_n), .Y(N101) );
  INVX1 U13600 ( .A(tmp_7_reg_1544[30]), .Y(n10807) );
  INVX1 U13601 ( .A(tmp_7_reg_1544[26]), .Y(n10803) );
  INVX1 U13602 ( .A(tmp_7_reg_1544[22]), .Y(n10799) );
  INVX1 U13603 ( .A(tmp_7_reg_1544[18]), .Y(n10795) );
  INVX1 U13604 ( .A(tmp_7_reg_1544[14]), .Y(n10791) );
  INVX1 U13605 ( .A(tmp_7_reg_1544[10]), .Y(n10787) );
  INVX1 U13606 ( .A(tmp_7_reg_1544[6]), .Y(n10783) );
  INVX1 U13607 ( .A(tmp_7_reg_1544[2]), .Y(n10779) );
  INVX1 U13608 ( .A(tmp_6_reg_1538[30]), .Y(n10773) );
  INVX1 U13609 ( .A(tmp_6_reg_1538[26]), .Y(n10769) );
  INVX1 U13610 ( .A(tmp_6_reg_1538[22]), .Y(n10765) );
  INVX1 U13611 ( .A(tmp_6_reg_1538[18]), .Y(n10761) );
  INVX1 U13612 ( .A(tmp_6_reg_1538[14]), .Y(n10757) );
  INVX1 U13613 ( .A(tmp_6_reg_1538[10]), .Y(n10753) );
  INVX1 U13614 ( .A(tmp_6_reg_1538[6]), .Y(n10749) );
  INVX1 U13615 ( .A(tmp_6_reg_1538[2]), .Y(n10745) );
  INVX1 U13616 ( .A(tmp_7_reg_1544[4]), .Y(n10781) );
  INVX1 U13617 ( .A(tmp_6_reg_1538[4]), .Y(n10747) );
  INVX1 U13618 ( .A(recentdatapoints_len[0]), .Y(n9825) );
  INVX1 U13619 ( .A(recentABools_len[4]), .Y(n10608) );
  INVX1 U13620 ( .A(recentVBools_len[4]), .Y(n10113) );
  INVX1 U13621 ( .A(tmp_7_reg_1544[28]), .Y(n10805) );
  INVX1 U13622 ( .A(tmp_7_reg_1544[12]), .Y(n10789) );
  INVX1 U13623 ( .A(tmp_6_reg_1538[28]), .Y(n10771) );
  INVX1 U13624 ( .A(tmp_6_reg_1538[12]), .Y(n10755) );
  INVX1 U13625 ( .A(s_axi_AXILiteS_ARADDR[6]), .Y(n9317) );
  OR2X1 U13626 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[30]), .B(n8800), 
        .Y(n8844) );
  OR2X1 U13627 ( .A(CircularBuffer_sum_read_assign_reg_1610[30]), .B(n8807), 
        .Y(n8845) );
  INVX1 U13628 ( .A(tmp_7_reg_1544[20]), .Y(n10797) );
  INVX1 U13629 ( .A(tmp_7_reg_1544[16]), .Y(n10793) );
  INVX1 U13630 ( .A(tmp_6_reg_1538[20]), .Y(n10763) );
  INVX1 U13631 ( .A(tmp_6_reg_1538[16]), .Y(n10759) );
  INVX1 U13632 ( .A(tmp_7_reg_1544[21]), .Y(n10798) );
  INVX1 U13633 ( .A(tmp_7_reg_1544[17]), .Y(n10794) );
  INVX1 U13634 ( .A(tmp_7_reg_1544[5]), .Y(n10782) );
  INVX1 U13635 ( .A(tmp_6_reg_1538[21]), .Y(n10764) );
  INVX1 U13636 ( .A(tmp_6_reg_1538[17]), .Y(n10760) );
  INVX1 U13637 ( .A(tmp_6_reg_1538[5]), .Y(n10748) );
  INVX1 U13638 ( .A(recentABools_len[3]), .Y(n10607) );
  INVX1 U13639 ( .A(recentVBools_len[3]), .Y(n10112) );
  OR2X1 U13640 ( .A(AbeatDelay_new_reg_394[22]), .B(AbeatDelay_new_reg_394[21]), .Y(n11048) );
  OR2X1 U13641 ( .A(AbeatDelay_new_reg_394[22]), .B(AbeatDelay_new_reg_394[21]), .Y(n11068) );
  INVX1 U13642 ( .A(recentVBools_sum[31]), .Y(n10241) );
  AND2X1 U13643 ( .A(n11239), .B(n11238), .Y(n11240) );
  OR2X1 U13644 ( .A(p_tmp_i_reg_1556[9]), .B(p_tmp_i_reg_1556[8]), .Y(n11237)
         );
  INVX1 U13645 ( .A(\Decision_AXILiteS_s_axi_U/int_isr[1] ), .Y(n10884) );
  INVX1 U13646 ( .A(recentdatapoints_len[31]), .Y(n9858) );
  INVX1 U13647 ( .A(tmp_7_reg_1544[31]), .Y(n10808) );
  INVX1 U13648 ( .A(tmp_6_reg_1538[31]), .Y(n10774) );
  INVX1 U13649 ( .A(recentABools_len[31]), .Y(n10669) );
  INVX1 U13650 ( .A(recentVBools_len[31]), .Y(n10172) );
  INVX1 U13651 ( .A(tmp_38_i_reg_1550[4]), .Y(n9928) );
  INVX1 U13652 ( .A(recentABools_len[7]), .Y(n10611) );
  INVX1 U13653 ( .A(recentABools_len[18]), .Y(n10622) );
  INVX1 U13654 ( .A(recentVBools_len[7]), .Y(n10116) );
  INVX1 U13655 ( .A(recentVBools_len[18]), .Y(n10127) );
  INVX1 U13656 ( .A(recentdatapoints_len[7]), .Y(n9835) );
  INVX1 U13657 ( .A(tmp_7_reg_1544[9]), .Y(n10786) );
  INVX1 U13658 ( .A(tmp_6_reg_1538[9]), .Y(n10752) );
  INVX1 U13659 ( .A(tmp_7_reg_1544[29]), .Y(n10806) );
  INVX1 U13660 ( .A(tmp_7_reg_1544[25]), .Y(n10802) );
  INVX1 U13661 ( .A(tmp_7_reg_1544[13]), .Y(n10790) );
  INVX1 U13662 ( .A(tmp_6_reg_1538[29]), .Y(n10772) );
  INVX1 U13663 ( .A(tmp_6_reg_1538[25]), .Y(n10768) );
  INVX1 U13664 ( .A(tmp_6_reg_1538[13]), .Y(n10756) );
  OR2X1 U13665 ( .A(VbeatFallDelay_new_1_reg_342[30]), .B(
        VbeatFallDelay_new_1_reg_342[29]), .Y(n11900) );
  INVX1 U13666 ( .A(\toReturn_8_reg_1755[0] ), .Y(n9383) );
  INVX1 U13667 ( .A(recentABools_sum[31]), .Y(n9384) );
  INVX1 U13668 ( .A(recentABools_len[6]), .Y(n10610) );
  INVX1 U13669 ( .A(recentABools_len[17]), .Y(n10621) );
  INVX1 U13670 ( .A(recentVBools_len[6]), .Y(n10115) );
  INVX1 U13671 ( .A(recentVBools_len[17]), .Y(n10126) );
  INVX1 U13672 ( .A(recentdatapoints_len[6]), .Y(n9834) );
  OR2X1 U13673 ( .A(s_axi_AXILiteS_ARADDR[1]), .B(s_axi_AXILiteS_ARADDR[0]), 
        .Y(\Decision_AXILiteS_s_axi_U/n315 ) );
  INVX1 U13674 ( .A(tmp_38_i_reg_1550[2]), .Y(n9830) );
  INVX1 U13675 ( .A(\toReturn_7_reg_1750[0] ), .Y(n10667) );
  INVX1 U13676 ( .A(\toReturn_5_reg_1655[0] ), .Y(n10207) );
  INVX1 U13677 ( .A(\toReturn_6_reg_1660[0] ), .Y(n10205) );
  INVX1 U13678 ( .A(\recentABools_data_load_reg_1700[0] ), .Y(n10666) );
  INVX1 U13679 ( .A(\recentVBools_data_load_reg_1584[0] ), .Y(n10206) );
  INVX1 U13680 ( .A(recentABools_len[30]), .Y(n10573) );
  INVX1 U13681 ( .A(recentABools_len[5]), .Y(n10609) );
  INVX1 U13682 ( .A(recentABools_len[28]), .Y(n10632) );
  INVX1 U13683 ( .A(recentABools_len[24]), .Y(n10628) );
  INVX1 U13684 ( .A(recentABools_len[14]), .Y(n10618) );
  INVX1 U13685 ( .A(recentABools_len[16]), .Y(n10620) );
  INVX1 U13686 ( .A(recentABools_len[12]), .Y(n10616) );
  INVX1 U13687 ( .A(recentVBools_len[30]), .Y(n10078) );
  INVX1 U13688 ( .A(recentVBools_len[5]), .Y(n10114) );
  INVX1 U13689 ( .A(recentVBools_len[28]), .Y(n10137) );
  INVX1 U13690 ( .A(recentVBools_len[24]), .Y(n10133) );
  INVX1 U13691 ( .A(recentVBools_len[14]), .Y(n10123) );
  INVX1 U13692 ( .A(recentVBools_len[16]), .Y(n10125) );
  INVX1 U13693 ( .A(recentVBools_len[12]), .Y(n10121) );
  INVX1 U13694 ( .A(recentdatapoints_len[12]), .Y(n9839) );
  INVX1 U13695 ( .A(recentdatapoints_len[14]), .Y(n9841) );
  INVX1 U13696 ( .A(recentdatapoints_len[21]), .Y(n9848) );
  INVX1 U13697 ( .A(recentdatapoints_len[18]), .Y(n9845) );
  INVX1 U13698 ( .A(recentdatapoints_len[5]), .Y(n9833) );
  INVX1 U13699 ( .A(recentdatapoints_len[29]), .Y(n9856) );
  INVX1 U13700 ( .A(recentdatapoints_len[25]), .Y(n9852) );
  INVX1 U13701 ( .A(recentABools_len[29]), .Y(n10633) );
  INVX1 U13702 ( .A(recentABools_len[27]), .Y(n10631) );
  INVX1 U13703 ( .A(recentABools_len[23]), .Y(n10627) );
  INVX1 U13704 ( .A(recentABools_len[13]), .Y(n10617) );
  INVX1 U13705 ( .A(recentABools_len[15]), .Y(n10619) );
  INVX1 U13706 ( .A(recentABools_len[11]), .Y(n10615) );
  INVX1 U13707 ( .A(recentVBools_len[29]), .Y(n10138) );
  INVX1 U13708 ( .A(recentVBools_len[27]), .Y(n10136) );
  INVX1 U13709 ( .A(recentVBools_len[23]), .Y(n10132) );
  INVX1 U13710 ( .A(recentVBools_len[13]), .Y(n10122) );
  INVX1 U13711 ( .A(recentVBools_len[15]), .Y(n10124) );
  INVX1 U13712 ( .A(recentVBools_len[11]), .Y(n10120) );
  INVX1 U13713 ( .A(recentdatapoints_len[11]), .Y(n9838) );
  INVX1 U13714 ( .A(recentdatapoints_len[13]), .Y(n9840) );
  INVX1 U13715 ( .A(recentdatapoints_len[20]), .Y(n9847) );
  INVX1 U13716 ( .A(recentdatapoints_len[17]), .Y(n9844) );
  INVX1 U13717 ( .A(recentdatapoints_len[30]), .Y(n9857) );
  INVX1 U13718 ( .A(recentdatapoints_len[3]), .Y(n9831) );
  INVX1 U13719 ( .A(recentdatapoints_len[28]), .Y(n9855) );
  INVX1 U13720 ( .A(recentdatapoints_len[24]), .Y(n9851) );
  INVX1 U13721 ( .A(tmp_38_i_reg_1550[19]), .Y(n9913) );
  INVX1 U13722 ( .A(tmp_38_i_reg_1550[21]), .Y(n9911) );
  OR2X1 U13723 ( .A(p_tmp_i_reg_1556[15]), .B(p_tmp_i_reg_1556[14]), .Y(n11247) );
  INVX1 U13724 ( .A(tmp_38_i_reg_1550[30]), .Y(n9902) );
  INVX1 U13725 ( .A(a_thresh[21]), .Y(n9781) );
  INVX1 U13726 ( .A(v_thresh[21]), .Y(n9522) );
  INVX1 U13727 ( .A(\Decision_AXILiteS_s_axi_U/waddr[2] ), .Y(n10894) );
  INVX1 U13728 ( .A(a_thresh[27]), .Y(n9787) );
  INVX1 U13729 ( .A(v_thresh[27]), .Y(n9529) );
  INVX1 U13730 ( .A(CircularBuffer_len_write_assig_2_reg_1729[7]), .Y(n10641)
         );
  INVX1 U13731 ( .A(CircularBuffer_len_write_assig_reg_1634[7]), .Y(n10146) );
  INVX1 U13732 ( .A(tmp_7_reg_1544[0]), .Y(n10777) );
  INVX1 U13733 ( .A(tmp_6_reg_1538[0]), .Y(n10743) );
  INVX1 U13734 ( .A(a_thresh[6]), .Y(n9770) );
  INVX1 U13735 ( .A(a_thresh[2]), .Y(n9767) );
  INVX1 U13736 ( .A(a_thresh[10]), .Y(n9772) );
  INVX1 U13737 ( .A(a_thresh[14]), .Y(n9775) );
  INVX1 U13738 ( .A(v_thresh[6]), .Y(n9504) );
  INVX1 U13739 ( .A(v_thresh[2]), .Y(n9499) );
  INVX1 U13740 ( .A(v_thresh[10]), .Y(n9510) );
  INVX1 U13741 ( .A(v_thresh[14]), .Y(n9516) );
  INVX1 U13742 ( .A(a_thresh[4]), .Y(n9768) );
  INVX1 U13743 ( .A(v_thresh[4]), .Y(n9500) );
  INVX1 U13744 ( .A(\last_sample_is_V_V[0] ), .Y(n10240) );
  INVX1 U13745 ( .A(\Decision_AXILiteS_s_axi_U/int_ier[0] ), .Y(n10886) );
  INVX1 U13746 ( .A(tmp_38_i_reg_1550[29]), .Y(n9903) );
  INVX1 U13747 ( .A(\Decision_AXILiteS_s_axi_U/int_gie ), .Y(n10888) );
  INVX1 U13748 ( .A(tmp_38_i_reg_1550[13]), .Y(n9919) );
  INVX1 U13749 ( .A(tmp_38_i_reg_1550[0]), .Y(n9859) );
  INVX1 U13750 ( .A(tmp_38_i_reg_1550[28]), .Y(n9904) );
  INVX1 U13751 ( .A(tmp_38_i_reg_1550[24]), .Y(n9908) );
  INVX1 U13752 ( .A(a_thresh[12]), .Y(n9773) );
  INVX1 U13753 ( .A(v_thresh[12]), .Y(n9512) );
  AND2X1 U13754 ( .A(s_axi_AXILiteS_WDATA[0]), .B(s_axi_AXILiteS_WSTRB[0]), 
        .Y(\Decision_AXILiteS_s_axi_U/n621 ) );
  INVX1 U13755 ( .A(n11908), .Y(n10367) );
  INVX1 U13756 ( .A(tmp_38_i_reg_1550[18]), .Y(n9914) );
  INVX1 U13757 ( .A(tmp_38_i_reg_1550[6]), .Y(n9926) );
  INVX1 U13758 ( .A(CircularBuffer_len_write_assig_2_reg_1729[9]), .Y(n10643)
         );
  INVX1 U13759 ( .A(CircularBuffer_len_write_assig_reg_1634[9]), .Y(n10148) );
  INVX1 U13760 ( .A(CircularBuffer_len_write_assig_2_reg_1729[17]), .Y(n10651)
         );
  INVX1 U13761 ( .A(CircularBuffer_len_write_assig_2_reg_1729[20]), .Y(n10654)
         );
  INVX1 U13762 ( .A(CircularBuffer_len_write_assig_2_reg_1729[24]), .Y(n10658)
         );
  INVX1 U13763 ( .A(CircularBuffer_len_write_assig_2_reg_1729[28]), .Y(n10662)
         );
  INVX1 U13764 ( .A(CircularBuffer_len_write_assig_reg_1634[17]), .Y(n10156)
         );
  INVX1 U13765 ( .A(CircularBuffer_len_write_assig_reg_1634[20]), .Y(n10159)
         );
  INVX1 U13766 ( .A(CircularBuffer_len_write_assig_reg_1634[24]), .Y(n10163)
         );
  INVX1 U13767 ( .A(CircularBuffer_len_write_assig_reg_1634[28]), .Y(n10167)
         );
  INVX1 U13768 ( .A(tmp_38_i_reg_1550[9]), .Y(n9923) );
  INVX1 U13769 ( .A(tmp_38_i_reg_1550[26]), .Y(n9906) );
  INVX1 U13770 ( .A(tmp_38_i_reg_1550[11]), .Y(n9921) );
  INVX1 U13771 ( .A(tmp_38_i_reg_1550[14]), .Y(n9918) );
  INVX1 U13772 ( .A(ap_CS_fsm[13]), .Y(n10670) );
  INVX1 U13773 ( .A(a_thresh[22]), .Y(n9782) );
  INVX1 U13774 ( .A(a_thresh[19]), .Y(n9779) );
  INVX1 U13775 ( .A(v_thresh[22]), .Y(n9523) );
  INVX1 U13776 ( .A(v_thresh[19]), .Y(n9520) );
  INVX1 U13777 ( .A(\recentABools_data_q0[0] ), .Y(n11047) );
  INVX1 U13778 ( .A(\recentVBools_data_q0[0] ), .Y(n11046) );
  INVX1 U13779 ( .A(CircularBuffer_len_write_assig_2_reg_1729[8]), .Y(n10642)
         );
  INVX1 U13780 ( .A(CircularBuffer_len_write_assig_reg_1634[8]), .Y(n10147) );
  INVX1 U13781 ( .A(CircularBuffer_len_write_assig_2_reg_1729[16]), .Y(n10650)
         );
  INVX1 U13782 ( .A(CircularBuffer_len_write_assig_2_reg_1729[23]), .Y(n10657)
         );
  INVX1 U13783 ( .A(CircularBuffer_len_write_assig_2_reg_1729[27]), .Y(n10661)
         );
  INVX1 U13784 ( .A(CircularBuffer_len_write_assig_reg_1634[16]), .Y(n10155)
         );
  INVX1 U13785 ( .A(CircularBuffer_len_write_assig_reg_1634[23]), .Y(n10162)
         );
  INVX1 U13786 ( .A(CircularBuffer_len_write_assig_reg_1634[27]), .Y(n10166)
         );
  INVX1 U13787 ( .A(tmp_38_i_reg_1550[8]), .Y(n9924) );
  INVX1 U13788 ( .A(tmp_38_i_reg_1550[20]), .Y(n9912) );
  INVX1 U13789 ( .A(a_thresh[13]), .Y(n9774) );
  INVX1 U13790 ( .A(v_thresh[13]), .Y(n9513) );
  INVX1 U13791 ( .A(a_thresh[5]), .Y(n9769) );
  INVX1 U13792 ( .A(v_thresh[5]), .Y(n9501) );
  INVX1 U13793 ( .A(CircularBuffer_len_write_assig_2_reg_1729[15]), .Y(n10649)
         );
  INVX1 U13794 ( .A(CircularBuffer_len_write_assig_reg_1634[15]), .Y(n10154)
         );
  INVX1 U13795 ( .A(a_thresh[9]), .Y(n9771) );
  INVX1 U13796 ( .A(v_thresh[9]), .Y(n9507) );
  INVX1 U13797 ( .A(tmp_38_i_reg_1550[1]), .Y(n9828) );
  INVX1 U13798 ( .A(n11256), .Y(n10303) );
  INVX1 U13799 ( .A(n11360), .Y(n10021) );
  INVX1 U13800 ( .A(n11412), .Y(n10330) );
  INVX1 U13801 ( .A(n11308), .Y(n9989) );
  INVX1 U13802 ( .A(CircularBuffer_len_write_assig_2_reg_1729[14]), .Y(n10648)
         );
  INVX1 U13803 ( .A(CircularBuffer_len_write_assig_reg_1634[14]), .Y(n10153)
         );
  INVX1 U13804 ( .A(tmp_38_i_reg_1550[31]), .Y(n9901) );
  INVX1 U13805 ( .A(tmp_38_i_reg_1550[3]), .Y(n9929) );
  INVX1 U13806 ( .A(tmp_38_i_reg_1550[27]), .Y(n9905) );
  INVX1 U13807 ( .A(tmp_38_i_reg_1550[12]), .Y(n9920) );
  INVX1 U13808 ( .A(tmp_38_i_reg_1550[15]), .Y(n9917) );
  INVX1 U13809 ( .A(tmp_38_i_reg_1550[17]), .Y(n9915) );
  INVX1 U13810 ( .A(tmp_38_i_reg_1550[16]), .Y(n9916) );
  INVX1 U13811 ( .A(tmp_38_i_reg_1550[5]), .Y(n9927) );
  INVX1 U13812 ( .A(tmp_38_i_reg_1550[23]), .Y(n9909) );
  INVX1 U13813 ( .A(\Decision_AXILiteS_s_axi_U/n633 ), .Y(n9275) );
  INVX1 U13814 ( .A(\Decision_AXILiteS_s_axi_U/n643 ), .Y(n9276) );
  INVX1 U13815 ( .A(aflip[7]), .Y(n9495) );
  INVX1 U13816 ( .A(vflip[3]), .Y(n9543) );
  INVX1 U13817 ( .A(vflip[7]), .Y(n9547) );
  INVX1 U13818 ( .A(aflip[2]), .Y(n9792) );
  INVX1 U13819 ( .A(aflip[6]), .Y(n9494) );
  INVX1 U13820 ( .A(vflip[2]), .Y(n9542) );
  INVX1 U13821 ( .A(vflip[6]), .Y(n9546) );
  INVX1 U13822 ( .A(\Decision_AXILiteS_s_axi_U/wstate[1] ), .Y(n10900) );
  INVX1 U13823 ( .A(\Decision_AXILiteS_s_axi_U/wstate[0] ), .Y(n10901) );
  INVX1 U13824 ( .A(\Decision_AXILiteS_s_axi_U/waddr[1] ), .Y(n10893) );
  INVX1 U13825 ( .A(tmp_3_reg_1589[31]), .Y(n10740) );
  INVX1 U13826 ( .A(tmp_3_reg_1589[30]), .Y(n10738) );
  INVX1 U13827 ( .A(tmp_3_reg_1589[29]), .Y(n10736) );
  INVX1 U13828 ( .A(tmp_3_reg_1589[28]), .Y(n10734) );
  INVX1 U13829 ( .A(tmp_3_reg_1589[27]), .Y(n10732) );
  INVX1 U13830 ( .A(tmp_3_reg_1589[26]), .Y(n10730) );
  INVX1 U13831 ( .A(tmp_3_reg_1589[25]), .Y(n10728) );
  INVX1 U13832 ( .A(tmp_3_reg_1589[24]), .Y(n10726) );
  INVX1 U13833 ( .A(tmp_3_reg_1589[23]), .Y(n10724) );
  INVX1 U13834 ( .A(tmp_3_reg_1589[22]), .Y(n10722) );
  INVX1 U13835 ( .A(tmp_3_reg_1589[21]), .Y(n10720) );
  INVX1 U13836 ( .A(tmp_3_reg_1589[20]), .Y(n10718) );
  INVX1 U13837 ( .A(tmp_3_reg_1589[19]), .Y(n10716) );
  INVX1 U13838 ( .A(tmp_3_reg_1589[18]), .Y(n10714) );
  INVX1 U13839 ( .A(tmp_3_reg_1589[17]), .Y(n10712) );
  INVX1 U13840 ( .A(tmp_3_reg_1589[16]), .Y(n10710) );
  INVX1 U13841 ( .A(tmp_3_reg_1589[15]), .Y(n10708) );
  INVX1 U13842 ( .A(tmp_3_reg_1589[14]), .Y(n10706) );
  INVX1 U13843 ( .A(tmp_3_reg_1589[13]), .Y(n10704) );
  INVX1 U13844 ( .A(tmp_3_reg_1589[12]), .Y(n10702) );
  INVX1 U13845 ( .A(tmp_3_reg_1589[11]), .Y(n10700) );
  INVX1 U13846 ( .A(tmp_3_reg_1589[10]), .Y(n10698) );
  INVX1 U13847 ( .A(tmp_3_reg_1589[9]), .Y(n10696) );
  INVX1 U13848 ( .A(tmp_3_reg_1589[8]), .Y(n10694) );
  INVX1 U13849 ( .A(tmp_3_reg_1589[7]), .Y(n10692) );
  INVX1 U13850 ( .A(tmp_3_reg_1589[6]), .Y(n10690) );
  INVX1 U13851 ( .A(tmp_3_reg_1589[5]), .Y(n10687) );
  INVX1 U13852 ( .A(tmp_3_reg_1589[4]), .Y(n10684) );
  INVX1 U13853 ( .A(tmp_3_reg_1589[3]), .Y(n10682) );
  INVX1 U13854 ( .A(tmp_3_reg_1589[2]), .Y(n10680) );
  INVX1 U13855 ( .A(tmp_3_reg_1589[1]), .Y(n10678) );
  INVX1 U13856 ( .A(tmp_3_reg_1589[0]), .Y(n10672) );
  INVX1 U13857 ( .A(tmp_4_reg_1596[31]), .Y(n10532) );
  INVX1 U13858 ( .A(tmp_4_reg_1596[30]), .Y(n10528) );
  INVX1 U13859 ( .A(tmp_4_reg_1596[29]), .Y(n10526) );
  INVX1 U13860 ( .A(tmp_4_reg_1596[28]), .Y(n10524) );
  INVX1 U13861 ( .A(tmp_4_reg_1596[27]), .Y(n10522) );
  INVX1 U13862 ( .A(tmp_4_reg_1596[26]), .Y(n10518) );
  INVX1 U13863 ( .A(tmp_4_reg_1596[25]), .Y(n10516) );
  INVX1 U13864 ( .A(tmp_4_reg_1596[24]), .Y(n10513) );
  INVX1 U13865 ( .A(tmp_4_reg_1596[23]), .Y(n10511) );
  INVX1 U13866 ( .A(tmp_4_reg_1596[22]), .Y(n10507) );
  INVX1 U13867 ( .A(tmp_4_reg_1596[21]), .Y(n10505) );
  INVX1 U13868 ( .A(tmp_4_reg_1596[20]), .Y(n10502) );
  INVX1 U13869 ( .A(tmp_4_reg_1596[19]), .Y(n10500) );
  INVX1 U13870 ( .A(tmp_4_reg_1596[18]), .Y(n10496) );
  INVX1 U13871 ( .A(tmp_4_reg_1596[17]), .Y(n10494) );
  INVX1 U13872 ( .A(tmp_4_reg_1596[16]), .Y(n10492) );
  INVX1 U13873 ( .A(tmp_4_reg_1596[15]), .Y(n10490) );
  INVX1 U13874 ( .A(tmp_4_reg_1596[14]), .Y(n10486) );
  INVX1 U13875 ( .A(tmp_4_reg_1596[13]), .Y(n10484) );
  INVX1 U13876 ( .A(tmp_4_reg_1596[12]), .Y(n10481) );
  INVX1 U13877 ( .A(tmp_4_reg_1596[11]), .Y(n10479) );
  INVX1 U13878 ( .A(tmp_4_reg_1596[10]), .Y(n10475) );
  INVX1 U13879 ( .A(tmp_4_reg_1596[9]), .Y(n10473) );
  INVX1 U13880 ( .A(tmp_4_reg_1596[8]), .Y(n10469) );
  INVX1 U13881 ( .A(tmp_4_reg_1596[7]), .Y(n10467) );
  INVX1 U13882 ( .A(tmp_4_reg_1596[6]), .Y(n10464) );
  INVX1 U13883 ( .A(tmp_4_reg_1596[5]), .Y(n10462) );
  INVX1 U13884 ( .A(tmp_4_reg_1596[4]), .Y(n10460) );
  INVX1 U13885 ( .A(tmp_4_reg_1596[3]), .Y(n10458) );
  INVX1 U13886 ( .A(tmp_4_reg_1596[2]), .Y(n10455) );
  INVX1 U13887 ( .A(tmp_4_reg_1596[1]), .Y(n10453) );
  INVX1 U13888 ( .A(tmp_4_reg_1596[0]), .Y(n10450) );
  INVX1 U13889 ( .A(tmp_5_reg_1603[31]), .Y(n10448) );
  INVX1 U13890 ( .A(tmp_5_reg_1603[30]), .Y(n10444) );
  INVX1 U13891 ( .A(tmp_5_reg_1603[29]), .Y(n10442) );
  INVX1 U13892 ( .A(tmp_5_reg_1603[28]), .Y(n10440) );
  INVX1 U13893 ( .A(tmp_5_reg_1603[27]), .Y(n10438) );
  INVX1 U13894 ( .A(tmp_5_reg_1603[26]), .Y(n10434) );
  INVX1 U13895 ( .A(tmp_5_reg_1603[25]), .Y(n10432) );
  INVX1 U13896 ( .A(tmp_5_reg_1603[24]), .Y(n10429) );
  INVX1 U13897 ( .A(tmp_5_reg_1603[23]), .Y(n10427) );
  INVX1 U13898 ( .A(tmp_5_reg_1603[22]), .Y(n10423) );
  INVX1 U13899 ( .A(tmp_5_reg_1603[21]), .Y(n10421) );
  INVX1 U13900 ( .A(tmp_5_reg_1603[20]), .Y(n10418) );
  INVX1 U13901 ( .A(tmp_5_reg_1603[19]), .Y(n10416) );
  INVX1 U13902 ( .A(tmp_5_reg_1603[18]), .Y(n10412) );
  INVX1 U13903 ( .A(tmp_5_reg_1603[17]), .Y(n10410) );
  INVX1 U13904 ( .A(tmp_5_reg_1603[16]), .Y(n10408) );
  INVX1 U13905 ( .A(tmp_5_reg_1603[15]), .Y(n10406) );
  INVX1 U13906 ( .A(tmp_5_reg_1603[14]), .Y(n10402) );
  INVX1 U13907 ( .A(tmp_5_reg_1603[13]), .Y(n10400) );
  INVX1 U13908 ( .A(tmp_5_reg_1603[12]), .Y(n10397) );
  INVX1 U13909 ( .A(tmp_5_reg_1603[11]), .Y(n10395) );
  INVX1 U13910 ( .A(tmp_5_reg_1603[10]), .Y(n10391) );
  INVX1 U13911 ( .A(tmp_5_reg_1603[9]), .Y(n10389) );
  INVX1 U13912 ( .A(tmp_5_reg_1603[8]), .Y(n10385) );
  INVX1 U13913 ( .A(tmp_5_reg_1603[7]), .Y(n10383) );
  INVX1 U13914 ( .A(tmp_5_reg_1603[6]), .Y(n10380) );
  INVX1 U13915 ( .A(tmp_5_reg_1603[5]), .Y(n10378) );
  INVX1 U13916 ( .A(tmp_5_reg_1603[4]), .Y(n10376) );
  INVX1 U13917 ( .A(tmp_5_reg_1603[3]), .Y(n10374) );
  INVX1 U13918 ( .A(tmp_5_reg_1603[2]), .Y(n10371) );
  INVX1 U13919 ( .A(tmp_5_reg_1603[1]), .Y(n10369) );
  INVX1 U13920 ( .A(tmp_5_reg_1603[0]), .Y(n10366) );
  INVX1 U13921 ( .A(aflip[3]), .Y(n9491) );
  INVX1 U13922 ( .A(\tmp_19_reg_409[0] ), .Y(n9385) );
  INVX1 U13923 ( .A(\Decision_AXILiteS_s_axi_U/rstate[0] ), .Y(
        s_axi_AXILiteS_ARREADY) );
  INVX1 U13924 ( .A(\Decision_AXILiteS_s_axi_U/waddr[0] ), .Y(n10892) );
  AND2X1 U13925 ( .A(ap_CS_fsm[10]), .B(ap_rst_n), .Y(N109) );
  AND2X1 U13926 ( .A(ap_CS_fsm[8]), .B(ap_rst_n), .Y(N107) );
  AND2X1 U13927 ( .A(ap_CS_fsm[5]), .B(ap_rst_n), .Y(N104) );
  AND2X1 U13928 ( .A(ap_CS_fsm[3]), .B(ap_rst_n), .Y(N102) );
  INVX1 U13929 ( .A(n11305), .Y(n10280) );
  INVX1 U13930 ( .A(n11409), .Y(n9998) );
  INVX1 U13931 ( .A(n11461), .Y(n10307) );
  INVX1 U13932 ( .A(n11357), .Y(n9966) );
  XNOR2X1 U13933 ( .A(n8591), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[10] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[10]) );
  XNOR2X1 U13934 ( .A(n8593), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[11] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[11]) );
  XNOR2X1 U13935 ( .A(n8595), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[12] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[12]) );
  XNOR2X1 U13936 ( .A(n8597), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[13] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[13]) );
  XNOR2X1 U13937 ( .A(n8599), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[14] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[14]) );
  XNOR2X1 U13938 ( .A(n8601), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[15] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[15]) );
  XNOR2X1 U13939 ( .A(n8603), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[16] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[16]) );
  XNOR2X1 U13940 ( .A(n8605), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[17] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[17]) );
  XNOR2X1 U13941 ( .A(n8607), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[18] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[18]) );
  XNOR2X1 U13942 ( .A(n8609), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[19] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[19]) );
  XNOR2X1 U13943 ( .A(n8576), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[1] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[1]) );
  XNOR2X1 U13944 ( .A(n8611), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[20] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[20]) );
  XNOR2X1 U13945 ( .A(n8613), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[21] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[21]) );
  XNOR2X1 U13946 ( .A(n8615), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[22] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[22]) );
  XNOR2X1 U13947 ( .A(n8617), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[23] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[23]) );
  XNOR2X1 U13948 ( .A(n8619), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[24] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[24]) );
  XNOR2X1 U13949 ( .A(n8621), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[25] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[25]) );
  XNOR2X1 U13950 ( .A(n8623), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[26] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[26]) );
  XNOR2X1 U13951 ( .A(n8625), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[27] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[27]) );
  XNOR2X1 U13952 ( .A(n8627), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[28] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[28]) );
  XNOR2X1 U13953 ( .A(n8629), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[29] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[29]) );
  XNOR2X1 U13954 ( .A(n8635), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[2] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[2]) );
  XNOR2X1 U13955 ( .A(n8631), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[30] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[30]) );
  XNOR2X1 U13956 ( .A(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[31] ), .B(
        n8846), .Y(CircularBuffer_sum_write_assig_3_fu_1242_p2[31]) );
  XNOR2X1 U13957 ( .A(n8578), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[3] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[3]) );
  XNOR2X1 U13958 ( .A(n8580), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[4] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[4]) );
  XNOR2X1 U13959 ( .A(n8581), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[5] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[5]) );
  XNOR2X1 U13960 ( .A(n8583), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[6] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[6]) );
  XNOR2X1 U13961 ( .A(n8585), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[7] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[7]) );
  XNOR2X1 U13962 ( .A(n8587), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[8] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[8]) );
  XNOR2X1 U13963 ( .A(n8589), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[9] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[9]) );
  XNOR2X1 U13964 ( .A(n9383), .B(
        \dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[0] ), .Y(
        CircularBuffer_sum_write_assig_3_fu_1242_p2[0]) );
  XNOR2X1 U13965 ( .A(n8688), .B(CircularBuffer_sum_read_assign_1_reg_1705[10]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[10] ) );
  XNOR2X1 U13966 ( .A(n8692), .B(CircularBuffer_sum_read_assign_1_reg_1705[11]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[11] ) );
  XNOR2X1 U13967 ( .A(n8696), .B(CircularBuffer_sum_read_assign_1_reg_1705[12]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[12] ) );
  XNOR2X1 U13968 ( .A(n8700), .B(CircularBuffer_sum_read_assign_1_reg_1705[13]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[13] ) );
  XNOR2X1 U13969 ( .A(n8704), .B(CircularBuffer_sum_read_assign_1_reg_1705[14]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[14] ) );
  XNOR2X1 U13970 ( .A(n8710), .B(CircularBuffer_sum_read_assign_1_reg_1705[15]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[15] ) );
  XNOR2X1 U13971 ( .A(n8716), .B(CircularBuffer_sum_read_assign_1_reg_1705[16]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[16] ) );
  XNOR2X1 U13972 ( .A(n8722), .B(CircularBuffer_sum_read_assign_1_reg_1705[17]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[17] ) );
  XNOR2X1 U13973 ( .A(n8728), .B(CircularBuffer_sum_read_assign_1_reg_1705[18]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[18] ) );
  XNOR2X1 U13974 ( .A(n8734), .B(CircularBuffer_sum_read_assign_1_reg_1705[19]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[19] ) );
  XNOR2X1 U13975 ( .A(n8667), .B(CircularBuffer_sum_read_assign_1_reg_1705[1]), 
        .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[1] ) );
  XNOR2X1 U13976 ( .A(n8740), .B(CircularBuffer_sum_read_assign_1_reg_1705[20]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[20] ) );
  XNOR2X1 U13977 ( .A(n8746), .B(CircularBuffer_sum_read_assign_1_reg_1705[21]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[21] ) );
  XNOR2X1 U13978 ( .A(n8752), .B(CircularBuffer_sum_read_assign_1_reg_1705[22]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[22] ) );
  XNOR2X1 U13979 ( .A(n8758), .B(CircularBuffer_sum_read_assign_1_reg_1705[23]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[23] ) );
  XNOR2X1 U13980 ( .A(n8764), .B(CircularBuffer_sum_read_assign_1_reg_1705[24]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[24] ) );
  XNOR2X1 U13981 ( .A(n8770), .B(CircularBuffer_sum_read_assign_1_reg_1705[25]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[25] ) );
  XNOR2X1 U13982 ( .A(n8776), .B(CircularBuffer_sum_read_assign_1_reg_1705[26]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[26] ) );
  XNOR2X1 U13983 ( .A(n8782), .B(CircularBuffer_sum_read_assign_1_reg_1705[27]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[27] ) );
  XNOR2X1 U13984 ( .A(n8788), .B(CircularBuffer_sum_read_assign_1_reg_1705[28]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[28] ) );
  XNOR2X1 U13985 ( .A(n8794), .B(CircularBuffer_sum_read_assign_1_reg_1705[29]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[29] ) );
  XNOR2X1 U13986 ( .A(n8837), .B(CircularBuffer_sum_read_assign_1_reg_1705[2]), 
        .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[2] ) );
  XNOR2X1 U13987 ( .A(n8800), .B(CircularBuffer_sum_read_assign_1_reg_1705[30]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[30] ) );
  XNOR2X1 U13988 ( .A(CircularBuffer_sum_read_assign_1_reg_1705[31]), .B(n8844), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[31] ) );
  XNOR2X1 U13989 ( .A(n8673), .B(CircularBuffer_sum_read_assign_1_reg_1705[3]), 
        .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[3] ) );
  XNOR2X1 U13990 ( .A(n8675), .B(CircularBuffer_sum_read_assign_1_reg_1705[4]), 
        .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[4] ) );
  XNOR2X1 U13991 ( .A(n8676), .B(CircularBuffer_sum_read_assign_1_reg_1705[5]), 
        .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[5] ) );
  XNOR2X1 U13992 ( .A(n8678), .B(CircularBuffer_sum_read_assign_1_reg_1705[6]), 
        .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[6] ) );
  XNOR2X1 U13993 ( .A(n8680), .B(CircularBuffer_sum_read_assign_1_reg_1705[7]), 
        .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[7] ) );
  XNOR2X1 U13994 ( .A(n8682), .B(CircularBuffer_sum_read_assign_1_reg_1705[8]), 
        .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[8] ) );
  XNOR2X1 U13995 ( .A(n8684), .B(CircularBuffer_sum_read_assign_1_reg_1705[9]), 
        .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[9] ) );
  XNOR2X1 U13996 ( .A(n10667), .B(CircularBuffer_sum_read_assign_1_reg_1705[0]), .Y(\dp_cluster_3/CircularBuffer_sum_write_assig_2_fu_1234_p2[0] ) );
  XNOR2X1 U13997 ( .A(n8594), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[10] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[10]) );
  XNOR2X1 U13998 ( .A(n8596), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[11] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[11]) );
  XNOR2X1 U13999 ( .A(n8598), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[12] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[12]) );
  XNOR2X1 U14000 ( .A(n8600), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[13] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[13]) );
  XNOR2X1 U14001 ( .A(n8602), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[14] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[14]) );
  XNOR2X1 U14002 ( .A(n8604), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[15] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[15]) );
  XNOR2X1 U14003 ( .A(n8606), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[16] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[16]) );
  XNOR2X1 U14004 ( .A(n8608), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[17] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[17]) );
  XNOR2X1 U14005 ( .A(n8610), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[18] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[18]) );
  XNOR2X1 U14006 ( .A(n8612), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[19] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[19]) );
  XNOR2X1 U14007 ( .A(n8577), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[1] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[1]) );
  XNOR2X1 U14008 ( .A(n8614), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[20] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[20]) );
  XNOR2X1 U14009 ( .A(n8616), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[21] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[21]) );
  XNOR2X1 U14010 ( .A(n8618), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[22] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[22]) );
  XNOR2X1 U14011 ( .A(n8620), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[23] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[23]) );
  XNOR2X1 U14012 ( .A(n8622), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[24] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[24]) );
  XNOR2X1 U14013 ( .A(n8624), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[25] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[25]) );
  XNOR2X1 U14014 ( .A(n8626), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[26] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[26]) );
  XNOR2X1 U14015 ( .A(n8628), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[27] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[27]) );
  XNOR2X1 U14016 ( .A(n8630), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[28] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[28]) );
  XNOR2X1 U14017 ( .A(n8632), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[29] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[29]) );
  XNOR2X1 U14018 ( .A(n8634), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[2] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[2]) );
  XNOR2X1 U14019 ( .A(n8633), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[30] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[30]) );
  XNOR2X1 U14020 ( .A(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[31] ), .B(n8847), .Y(CircularBuffer_sum_write_assig_1_fu_917_p2[31]) );
  XNOR2X1 U14021 ( .A(n8579), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[3] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[3]) );
  XNOR2X1 U14022 ( .A(n8582), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[4] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[4]) );
  XNOR2X1 U14023 ( .A(n8584), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[5] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[5]) );
  XNOR2X1 U14024 ( .A(n8586), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[6] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[6]) );
  XNOR2X1 U14025 ( .A(n8588), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[7] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[7]) );
  XNOR2X1 U14026 ( .A(n8590), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[8] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[8]) );
  XNOR2X1 U14027 ( .A(n8592), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[9] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[9]) );
  XNOR2X1 U14028 ( .A(n10205), .B(
        \dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[0] ), .Y(
        CircularBuffer_sum_write_assig_1_fu_917_p2[0]) );
  XNOR2X1 U14029 ( .A(n8693), .B(CircularBuffer_sum_read_assign_reg_1610[10]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[10] ) );
  XNOR2X1 U14030 ( .A(n8697), .B(CircularBuffer_sum_read_assign_reg_1610[11]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[11] ) );
  XNOR2X1 U14031 ( .A(n8701), .B(CircularBuffer_sum_read_assign_reg_1610[12]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[12] ) );
  XNOR2X1 U14032 ( .A(n8706), .B(CircularBuffer_sum_read_assign_reg_1610[13]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[13] ) );
  XNOR2X1 U14033 ( .A(n8712), .B(CircularBuffer_sum_read_assign_reg_1610[14]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[14] ) );
  XNOR2X1 U14034 ( .A(n8718), .B(CircularBuffer_sum_read_assign_reg_1610[15]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[15] ) );
  XNOR2X1 U14035 ( .A(n8724), .B(CircularBuffer_sum_read_assign_reg_1610[16]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[16] ) );
  XNOR2X1 U14036 ( .A(n8730), .B(CircularBuffer_sum_read_assign_reg_1610[17]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[17] ) );
  XNOR2X1 U14037 ( .A(n8736), .B(CircularBuffer_sum_read_assign_reg_1610[18]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[18] ) );
  XNOR2X1 U14038 ( .A(n8742), .B(CircularBuffer_sum_read_assign_reg_1610[19]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[19] ) );
  XNOR2X1 U14039 ( .A(n8668), .B(CircularBuffer_sum_read_assign_reg_1610[1]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[1] ) );
  XNOR2X1 U14040 ( .A(n8748), .B(CircularBuffer_sum_read_assign_reg_1610[20]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[20] ) );
  XNOR2X1 U14041 ( .A(n8754), .B(CircularBuffer_sum_read_assign_reg_1610[21]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[21] ) );
  XNOR2X1 U14042 ( .A(n8760), .B(CircularBuffer_sum_read_assign_reg_1610[22]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[22] ) );
  XNOR2X1 U14043 ( .A(n8766), .B(CircularBuffer_sum_read_assign_reg_1610[23]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[23] ) );
  XNOR2X1 U14044 ( .A(n8772), .B(CircularBuffer_sum_read_assign_reg_1610[24]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[24] ) );
  XNOR2X1 U14045 ( .A(n8778), .B(CircularBuffer_sum_read_assign_reg_1610[25]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[25] ) );
  XNOR2X1 U14046 ( .A(n8784), .B(CircularBuffer_sum_read_assign_reg_1610[26]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[26] ) );
  XNOR2X1 U14047 ( .A(n8790), .B(CircularBuffer_sum_read_assign_reg_1610[27]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[27] ) );
  XNOR2X1 U14048 ( .A(n8796), .B(CircularBuffer_sum_read_assign_reg_1610[28]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[28] ) );
  XNOR2X1 U14049 ( .A(n8802), .B(CircularBuffer_sum_read_assign_reg_1610[29]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[29] ) );
  XNOR2X1 U14050 ( .A(n8838), .B(CircularBuffer_sum_read_assign_reg_1610[2]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[2] ) );
  XNOR2X1 U14051 ( .A(n8807), .B(CircularBuffer_sum_read_assign_reg_1610[30]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[30] ) );
  XNOR2X1 U14052 ( .A(CircularBuffer_sum_read_assign_reg_1610[31]), .B(n8845), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[31] ) );
  XNOR2X1 U14053 ( .A(n8674), .B(CircularBuffer_sum_read_assign_reg_1610[3]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[3] ) );
  XNOR2X1 U14054 ( .A(n8677), .B(CircularBuffer_sum_read_assign_reg_1610[4]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[4] ) );
  XNOR2X1 U14055 ( .A(n8679), .B(CircularBuffer_sum_read_assign_reg_1610[5]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[5] ) );
  XNOR2X1 U14056 ( .A(n8681), .B(CircularBuffer_sum_read_assign_reg_1610[6]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[6] ) );
  XNOR2X1 U14057 ( .A(n8683), .B(CircularBuffer_sum_read_assign_reg_1610[7]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[7] ) );
  XNOR2X1 U14058 ( .A(n8685), .B(CircularBuffer_sum_read_assign_reg_1610[8]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[8] ) );
  XNOR2X1 U14059 ( .A(n8689), .B(CircularBuffer_sum_read_assign_reg_1610[9]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[9] ) );
  XNOR2X1 U14060 ( .A(n10207), .B(CircularBuffer_sum_read_assign_reg_1610[0]), 
        .Y(\dp_cluster_2/CircularBuffer_sum_write_assig_fu_909_p2[0] ) );
  XNOR2X1 U14061 ( .A(i_8_fu_1148_p2[1]), .B(i_8_fu_1148_p2[2]), .Y(
        i_9_fu_1160_p2[2]) );
  XNOR2X1 U14062 ( .A(n8638), .B(i_8_fu_1148_p2[3]), .Y(i_9_fu_1160_p2[3]) );
  XNOR2X1 U14063 ( .A(i_8_fu_1148_p2[4]), .B(n8642), .Y(i_9_fu_1160_p2[4]) );
  XNOR2X1 U14064 ( .A(n10541), .B(CircularBuffer_head_i_read_ass_1_reg_1719[0]), .Y(i_9_fu_1160_p2[0]) );
  XNOR2X1 U14065 ( .A(i_5_fu_854_p2[1]), .B(i_5_fu_854_p2[2]), .Y(
        i_6_fu_866_p2[2]) );
  XNOR2X1 U14066 ( .A(n8641), .B(i_5_fu_854_p2[3]), .Y(i_6_fu_866_p2[3]) );
  XNOR2X1 U14067 ( .A(i_5_fu_854_p2[4]), .B(n8848), .Y(i_6_fu_866_p2[4]) );
  XNOR2X1 U14068 ( .A(n10139), .B(CircularBuffer_head_i_read_ass_reg_1624[0]), 
        .Y(i_6_fu_866_p2[0]) );
  XNOR2X1 U14069 ( .A(i_2_fu_823_p2[1]), .B(i_2_fu_823_p2[2]), .Y(
        i_3_fu_835_p2[2]) );
  XNOR2X1 U14070 ( .A(n8639), .B(i_2_fu_823_p2[3]), .Y(i_3_fu_835_p2[3]) );
  XNOR2X1 U14071 ( .A(i_2_fu_823_p2[4]), .B(n8643), .Y(i_3_fu_835_p2[4]) );
  XNOR2X1 U14072 ( .A(n10076), .B(CircularBuffer_head_i_read_ass_reg_1624[0]), 
        .Y(i_3_fu_835_p2[0]) );
  XNOR2X1 U14073 ( .A(i_11_fu_1179_p2[1]), .B(i_11_fu_1179_p2[2]), .Y(
        i_12_fu_1191_p2[2]) );
  XNOR2X1 U14074 ( .A(n8640), .B(i_11_fu_1179_p2[3]), .Y(i_12_fu_1191_p2[3])
         );
  XNOR2X1 U14075 ( .A(i_11_fu_1179_p2[4]), .B(n8849), .Y(i_12_fu_1191_p2[4])
         );
  XNOR2X1 U14076 ( .A(n10634), .B(CircularBuffer_head_i_read_ass_1_reg_1719[0]), .Y(i_12_fu_1191_p2[0]) );
  XNOR2X1 U14077 ( .A(p_tmp_i_reg_1556[0]), .B(p_tmp_i_reg_1556[1]), .Y(
        i_1_fu_620_p2[1]) );
  XNOR2X1 U14078 ( .A(p_tmp_i_reg_1556[4]), .B(n8854), .Y(i_1_fu_620_p2[4]) );
  XNOR2X1 U14079 ( .A(n8721), .B(recentVBools_sum[10]), .Y(
        tmp_29_i_fu_752_p2[10]) );
  XNOR2X1 U14080 ( .A(n8727), .B(recentVBools_sum[11]), .Y(
        tmp_29_i_fu_752_p2[11]) );
  XNOR2X1 U14081 ( .A(n8733), .B(recentVBools_sum[12]), .Y(
        tmp_29_i_fu_752_p2[12]) );
  XNOR2X1 U14082 ( .A(n8739), .B(recentVBools_sum[13]), .Y(
        tmp_29_i_fu_752_p2[13]) );
  XNOR2X1 U14083 ( .A(n8745), .B(recentVBools_sum[14]), .Y(
        tmp_29_i_fu_752_p2[14]) );
  XNOR2X1 U14084 ( .A(n8751), .B(recentVBools_sum[15]), .Y(
        tmp_29_i_fu_752_p2[15]) );
  XNOR2X1 U14085 ( .A(n8757), .B(recentVBools_sum[16]), .Y(
        tmp_29_i_fu_752_p2[16]) );
  XNOR2X1 U14086 ( .A(n8763), .B(recentVBools_sum[17]), .Y(
        tmp_29_i_fu_752_p2[17]) );
  XNOR2X1 U14087 ( .A(n8769), .B(recentVBools_sum[18]), .Y(
        tmp_29_i_fu_752_p2[18]) );
  XNOR2X1 U14088 ( .A(n8775), .B(recentVBools_sum[19]), .Y(
        tmp_29_i_fu_752_p2[19]) );
  XNOR2X1 U14089 ( .A(n8670), .B(recentVBools_sum[1]), .Y(
        tmp_29_i_fu_752_p2[1]) );
  XNOR2X1 U14090 ( .A(n8781), .B(recentVBools_sum[20]), .Y(
        tmp_29_i_fu_752_p2[20]) );
  XNOR2X1 U14091 ( .A(n8787), .B(recentVBools_sum[21]), .Y(
        tmp_29_i_fu_752_p2[21]) );
  XNOR2X1 U14092 ( .A(n8793), .B(recentVBools_sum[22]), .Y(
        tmp_29_i_fu_752_p2[22]) );
  XNOR2X1 U14093 ( .A(n8799), .B(recentVBools_sum[23]), .Y(
        tmp_29_i_fu_752_p2[23]) );
  XNOR2X1 U14094 ( .A(n8805), .B(recentVBools_sum[24]), .Y(
        tmp_29_i_fu_752_p2[24]) );
  XNOR2X1 U14095 ( .A(n8810), .B(recentVBools_sum[25]), .Y(
        tmp_29_i_fu_752_p2[25]) );
  XNOR2X1 U14096 ( .A(n8814), .B(recentVBools_sum[26]), .Y(
        tmp_29_i_fu_752_p2[26]) );
  XNOR2X1 U14097 ( .A(n8818), .B(recentVBools_sum[27]), .Y(
        tmp_29_i_fu_752_p2[27]) );
  XNOR2X1 U14098 ( .A(n8822), .B(recentVBools_sum[28]), .Y(
        tmp_29_i_fu_752_p2[28]) );
  XNOR2X1 U14099 ( .A(n8826), .B(recentVBools_sum[29]), .Y(
        tmp_29_i_fu_752_p2[29]) );
  XNOR2X1 U14100 ( .A(n8840), .B(recentVBools_sum[2]), .Y(
        tmp_29_i_fu_752_p2[2]) );
  XNOR2X1 U14101 ( .A(n8830), .B(recentVBools_sum[30]), .Y(
        tmp_29_i_fu_752_p2[30]) );
  XNOR2X1 U14102 ( .A(recentVBools_sum[31]), .B(n8850), .Y(
        tmp_29_i_fu_752_p2[31]) );
  XNOR2X1 U14103 ( .A(n8687), .B(recentVBools_sum[3]), .Y(
        tmp_29_i_fu_752_p2[3]) );
  XNOR2X1 U14104 ( .A(n8691), .B(recentVBools_sum[4]), .Y(
        tmp_29_i_fu_752_p2[4]) );
  XNOR2X1 U14105 ( .A(n8695), .B(recentVBools_sum[5]), .Y(
        tmp_29_i_fu_752_p2[5]) );
  XNOR2X1 U14106 ( .A(n8699), .B(recentVBools_sum[6]), .Y(
        tmp_29_i_fu_752_p2[6]) );
  XNOR2X1 U14107 ( .A(n8703), .B(recentVBools_sum[7]), .Y(
        tmp_29_i_fu_752_p2[7]) );
  XNOR2X1 U14108 ( .A(n8709), .B(recentVBools_sum[8]), .Y(
        tmp_29_i_fu_752_p2[8]) );
  XNOR2X1 U14109 ( .A(n8715), .B(recentVBools_sum[9]), .Y(
        tmp_29_i_fu_752_p2[9]) );
  XNOR2X1 U14110 ( .A(n10206), .B(recentVBools_sum[0]), .Y(
        tmp_29_i_fu_752_p2[0]) );
  XNOR2X1 U14111 ( .A(n8720), .B(recentABools_sum[10]), .Y(
        tmp_29_i1_fu_1065_p2[10]) );
  XNOR2X1 U14112 ( .A(n8726), .B(recentABools_sum[11]), .Y(
        tmp_29_i1_fu_1065_p2[11]) );
  XNOR2X1 U14113 ( .A(n8732), .B(recentABools_sum[12]), .Y(
        tmp_29_i1_fu_1065_p2[12]) );
  XNOR2X1 U14114 ( .A(n8738), .B(recentABools_sum[13]), .Y(
        tmp_29_i1_fu_1065_p2[13]) );
  XNOR2X1 U14115 ( .A(n8744), .B(recentABools_sum[14]), .Y(
        tmp_29_i1_fu_1065_p2[14]) );
  XNOR2X1 U14116 ( .A(n8750), .B(recentABools_sum[15]), .Y(
        tmp_29_i1_fu_1065_p2[15]) );
  XNOR2X1 U14117 ( .A(n8756), .B(recentABools_sum[16]), .Y(
        tmp_29_i1_fu_1065_p2[16]) );
  XNOR2X1 U14118 ( .A(n8762), .B(recentABools_sum[17]), .Y(
        tmp_29_i1_fu_1065_p2[17]) );
  XNOR2X1 U14119 ( .A(n8768), .B(recentABools_sum[18]), .Y(
        tmp_29_i1_fu_1065_p2[18]) );
  XNOR2X1 U14120 ( .A(n8774), .B(recentABools_sum[19]), .Y(
        tmp_29_i1_fu_1065_p2[19]) );
  XNOR2X1 U14121 ( .A(n8669), .B(recentABools_sum[1]), .Y(
        tmp_29_i1_fu_1065_p2[1]) );
  XNOR2X1 U14122 ( .A(n8780), .B(recentABools_sum[20]), .Y(
        tmp_29_i1_fu_1065_p2[20]) );
  XNOR2X1 U14123 ( .A(n8786), .B(recentABools_sum[21]), .Y(
        tmp_29_i1_fu_1065_p2[21]) );
  XNOR2X1 U14124 ( .A(n8792), .B(recentABools_sum[22]), .Y(
        tmp_29_i1_fu_1065_p2[22]) );
  XNOR2X1 U14125 ( .A(n8798), .B(recentABools_sum[23]), .Y(
        tmp_29_i1_fu_1065_p2[23]) );
  XNOR2X1 U14126 ( .A(n8804), .B(recentABools_sum[24]), .Y(
        tmp_29_i1_fu_1065_p2[24]) );
  XNOR2X1 U14127 ( .A(n8809), .B(recentABools_sum[25]), .Y(
        tmp_29_i1_fu_1065_p2[25]) );
  XNOR2X1 U14128 ( .A(n8813), .B(recentABools_sum[26]), .Y(
        tmp_29_i1_fu_1065_p2[26]) );
  XNOR2X1 U14129 ( .A(n8817), .B(recentABools_sum[27]), .Y(
        tmp_29_i1_fu_1065_p2[27]) );
  XNOR2X1 U14130 ( .A(n8821), .B(recentABools_sum[28]), .Y(
        tmp_29_i1_fu_1065_p2[28]) );
  XNOR2X1 U14131 ( .A(n8825), .B(recentABools_sum[29]), .Y(
        tmp_29_i1_fu_1065_p2[29]) );
  XNOR2X1 U14132 ( .A(n8839), .B(recentABools_sum[2]), .Y(
        tmp_29_i1_fu_1065_p2[2]) );
  XNOR2X1 U14133 ( .A(n8829), .B(recentABools_sum[30]), .Y(
        tmp_29_i1_fu_1065_p2[30]) );
  XNOR2X1 U14134 ( .A(recentABools_sum[31]), .B(n8851), .Y(
        tmp_29_i1_fu_1065_p2[31]) );
  XNOR2X1 U14135 ( .A(n8686), .B(recentABools_sum[3]), .Y(
        tmp_29_i1_fu_1065_p2[3]) );
  XNOR2X1 U14136 ( .A(n8690), .B(recentABools_sum[4]), .Y(
        tmp_29_i1_fu_1065_p2[4]) );
  XNOR2X1 U14137 ( .A(n8694), .B(recentABools_sum[5]), .Y(
        tmp_29_i1_fu_1065_p2[5]) );
  XNOR2X1 U14138 ( .A(n8698), .B(recentABools_sum[6]), .Y(
        tmp_29_i1_fu_1065_p2[6]) );
  XNOR2X1 U14139 ( .A(n8702), .B(recentABools_sum[7]), .Y(
        tmp_29_i1_fu_1065_p2[7]) );
  XNOR2X1 U14140 ( .A(n8708), .B(recentABools_sum[8]), .Y(
        tmp_29_i1_fu_1065_p2[8]) );
  XNOR2X1 U14141 ( .A(n8714), .B(recentABools_sum[9]), .Y(
        tmp_29_i1_fu_1065_p2[9]) );
  XNOR2X1 U14142 ( .A(n10666), .B(recentABools_sum[0]), .Y(
        tmp_29_i1_fu_1065_p2[0]) );
  XNOR2X1 U14143 ( .A(CircularBuffer_len_read_assign_3_reg_1711[1]), .B(
        CircularBuffer_len_read_assign_3_reg_1711[2]), .Y(
        CircularBuffer_len_write_assig_3_fu_1249_p2[2]) );
  XNOR2X1 U14144 ( .A(n8841), .B(CircularBuffer_len_read_assign_3_reg_1711[3]), 
        .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[3]) );
  XNOR2X1 U14145 ( .A(n8671), .B(CircularBuffer_len_read_assign_3_reg_1711[4]), 
        .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[4]) );
  XNOR2X1 U14146 ( .A(n8835), .B(CircularBuffer_len_read_assign_3_reg_1711[5]), 
        .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[5]) );
  XNOR2X1 U14147 ( .A(n8705), .B(CircularBuffer_len_read_assign_3_reg_1711[6]), 
        .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[6]) );
  XNOR2X1 U14148 ( .A(n8711), .B(CircularBuffer_len_read_assign_3_reg_1711[7]), 
        .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[7]) );
  XNOR2X1 U14149 ( .A(n8717), .B(CircularBuffer_len_read_assign_3_reg_1711[8]), 
        .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[8]) );
  XNOR2X1 U14150 ( .A(n8723), .B(CircularBuffer_len_read_assign_3_reg_1711[9]), 
        .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[9]) );
  XNOR2X1 U14151 ( .A(n8729), .B(CircularBuffer_len_read_assign_3_reg_1711[10]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[10]) );
  XNOR2X1 U14152 ( .A(n8735), .B(CircularBuffer_len_read_assign_3_reg_1711[11]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[11]) );
  XNOR2X1 U14153 ( .A(n8741), .B(CircularBuffer_len_read_assign_3_reg_1711[12]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[12]) );
  XNOR2X1 U14154 ( .A(n8747), .B(CircularBuffer_len_read_assign_3_reg_1711[13]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[13]) );
  XNOR2X1 U14155 ( .A(n8753), .B(CircularBuffer_len_read_assign_3_reg_1711[14]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[14]) );
  XNOR2X1 U14156 ( .A(n8759), .B(CircularBuffer_len_read_assign_3_reg_1711[15]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[15]) );
  XNOR2X1 U14157 ( .A(n8765), .B(CircularBuffer_len_read_assign_3_reg_1711[16]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[16]) );
  XNOR2X1 U14158 ( .A(n8771), .B(CircularBuffer_len_read_assign_3_reg_1711[17]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[17]) );
  XNOR2X1 U14159 ( .A(n8777), .B(CircularBuffer_len_read_assign_3_reg_1711[18]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[18]) );
  XNOR2X1 U14160 ( .A(n8783), .B(CircularBuffer_len_read_assign_3_reg_1711[19]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[19]) );
  XNOR2X1 U14161 ( .A(n8789), .B(CircularBuffer_len_read_assign_3_reg_1711[20]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[20]) );
  XNOR2X1 U14162 ( .A(n8795), .B(CircularBuffer_len_read_assign_3_reg_1711[21]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[21]) );
  XNOR2X1 U14163 ( .A(n8801), .B(CircularBuffer_len_read_assign_3_reg_1711[22]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[22]) );
  XNOR2X1 U14164 ( .A(n8806), .B(CircularBuffer_len_read_assign_3_reg_1711[23]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[23]) );
  XNOR2X1 U14165 ( .A(n8811), .B(CircularBuffer_len_read_assign_3_reg_1711[24]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[24]) );
  XNOR2X1 U14166 ( .A(n8815), .B(CircularBuffer_len_read_assign_3_reg_1711[25]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[25]) );
  XNOR2X1 U14167 ( .A(n8819), .B(CircularBuffer_len_read_assign_3_reg_1711[26]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[26]) );
  XNOR2X1 U14168 ( .A(n8823), .B(CircularBuffer_len_read_assign_3_reg_1711[27]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[27]) );
  XNOR2X1 U14169 ( .A(n8827), .B(CircularBuffer_len_read_assign_3_reg_1711[28]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[28]) );
  XNOR2X1 U14170 ( .A(n8831), .B(CircularBuffer_len_read_assign_3_reg_1711[29]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[29]) );
  XNOR2X1 U14171 ( .A(n8833), .B(CircularBuffer_len_read_assign_3_reg_1711[30]), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[30]) );
  XNOR2X1 U14172 ( .A(CircularBuffer_len_read_assign_3_reg_1711[31]), .B(n8852), .Y(CircularBuffer_len_write_assig_3_fu_1249_p2[31]) );
  XNOR2X1 U14173 ( .A(CircularBuffer_len_read_assign_1_reg_1616[1]), .B(
        CircularBuffer_len_read_assign_1_reg_1616[2]), .Y(
        CircularBuffer_len_write_assig_1_fu_924_p2[2]) );
  XNOR2X1 U14174 ( .A(n8842), .B(CircularBuffer_len_read_assign_1_reg_1616[3]), 
        .Y(CircularBuffer_len_write_assig_1_fu_924_p2[3]) );
  XNOR2X1 U14175 ( .A(n8672), .B(CircularBuffer_len_read_assign_1_reg_1616[4]), 
        .Y(CircularBuffer_len_write_assig_1_fu_924_p2[4]) );
  XNOR2X1 U14176 ( .A(n8836), .B(CircularBuffer_len_read_assign_1_reg_1616[5]), 
        .Y(CircularBuffer_len_write_assig_1_fu_924_p2[5]) );
  XNOR2X1 U14177 ( .A(n8707), .B(CircularBuffer_len_read_assign_1_reg_1616[6]), 
        .Y(CircularBuffer_len_write_assig_1_fu_924_p2[6]) );
  XNOR2X1 U14178 ( .A(n8713), .B(CircularBuffer_len_read_assign_1_reg_1616[7]), 
        .Y(CircularBuffer_len_write_assig_1_fu_924_p2[7]) );
  XNOR2X1 U14179 ( .A(n8719), .B(CircularBuffer_len_read_assign_1_reg_1616[8]), 
        .Y(CircularBuffer_len_write_assig_1_fu_924_p2[8]) );
  XNOR2X1 U14180 ( .A(n8725), .B(CircularBuffer_len_read_assign_1_reg_1616[9]), 
        .Y(CircularBuffer_len_write_assig_1_fu_924_p2[9]) );
  XNOR2X1 U14181 ( .A(n8731), .B(CircularBuffer_len_read_assign_1_reg_1616[10]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[10]) );
  XNOR2X1 U14182 ( .A(n8737), .B(CircularBuffer_len_read_assign_1_reg_1616[11]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[11]) );
  XNOR2X1 U14183 ( .A(n8743), .B(CircularBuffer_len_read_assign_1_reg_1616[12]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[12]) );
  XNOR2X1 U14184 ( .A(n8749), .B(CircularBuffer_len_read_assign_1_reg_1616[13]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[13]) );
  XNOR2X1 U14185 ( .A(n8755), .B(CircularBuffer_len_read_assign_1_reg_1616[14]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[14]) );
  XNOR2X1 U14186 ( .A(n8761), .B(CircularBuffer_len_read_assign_1_reg_1616[15]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[15]) );
  XNOR2X1 U14187 ( .A(n8767), .B(CircularBuffer_len_read_assign_1_reg_1616[16]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[16]) );
  XNOR2X1 U14188 ( .A(n8773), .B(CircularBuffer_len_read_assign_1_reg_1616[17]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[17]) );
  XNOR2X1 U14189 ( .A(n8779), .B(CircularBuffer_len_read_assign_1_reg_1616[18]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[18]) );
  XNOR2X1 U14190 ( .A(n8785), .B(CircularBuffer_len_read_assign_1_reg_1616[19]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[19]) );
  XNOR2X1 U14191 ( .A(n8791), .B(CircularBuffer_len_read_assign_1_reg_1616[20]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[20]) );
  XNOR2X1 U14192 ( .A(n8797), .B(CircularBuffer_len_read_assign_1_reg_1616[21]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[21]) );
  XNOR2X1 U14193 ( .A(n8803), .B(CircularBuffer_len_read_assign_1_reg_1616[22]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[22]) );
  XNOR2X1 U14194 ( .A(n8808), .B(CircularBuffer_len_read_assign_1_reg_1616[23]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[23]) );
  XNOR2X1 U14195 ( .A(n8812), .B(CircularBuffer_len_read_assign_1_reg_1616[24]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[24]) );
  XNOR2X1 U14196 ( .A(n8816), .B(CircularBuffer_len_read_assign_1_reg_1616[25]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[25]) );
  XNOR2X1 U14197 ( .A(n8820), .B(CircularBuffer_len_read_assign_1_reg_1616[26]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[26]) );
  XNOR2X1 U14198 ( .A(n8824), .B(CircularBuffer_len_read_assign_1_reg_1616[27]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[27]) );
  XNOR2X1 U14199 ( .A(n8828), .B(CircularBuffer_len_read_assign_1_reg_1616[28]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[28]) );
  XNOR2X1 U14200 ( .A(n8832), .B(CircularBuffer_len_read_assign_1_reg_1616[29]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[29]) );
  XNOR2X1 U14201 ( .A(n8834), .B(CircularBuffer_len_read_assign_1_reg_1616[30]), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[30]) );
  XNOR2X1 U14202 ( .A(CircularBuffer_len_read_assign_1_reg_1616[31]), .B(n8853), .Y(CircularBuffer_len_write_assig_1_fu_924_p2[31]) );
  XOR2X1 U14203 ( .A(n8390), .B(n6944), .Y(datapointV_1_fu_674_p2[1]) );
  XOR2X1 U14204 ( .A(n8568), .B(n7261), .Y(datapointV_1_fu_674_p2[2]) );
  XOR2X1 U14205 ( .A(n8572), .B(n7638), .Y(datapointV_1_fu_674_p2[3]) );
  XOR2X1 U14206 ( .A(n8562), .B(n8101), .Y(datapointV_1_fu_674_p2[4]) );
  XOR2X1 U14207 ( .A(n8564), .B(n7857), .Y(datapointV_1_fu_674_p2[5]) );
  XOR2X1 U14208 ( .A(n8567), .B(n7435), .Y(datapointV_1_fu_674_p2[6]) );
  XOR2X1 U14209 ( .A(n8571), .B(n7096), .Y(datapointV_1_fu_674_p2[7]) );
  XOR2X1 U14210 ( .A(n8573), .B(n7436), .Y(datapointV_1_fu_674_p2[8]) );
  XOR2X1 U14211 ( .A(n8565), .B(n7856), .Y(datapointV_1_fu_674_p2[9]) );
  XOR2X1 U14212 ( .A(n8569), .B(n7097), .Y(datapointV_1_fu_674_p2[10]) );
  XOR2X1 U14213 ( .A(n8574), .B(n7262), .Y(datapointV_1_fu_674_p2[11]) );
  XOR2X1 U14214 ( .A(n8563), .B(n8387), .Y(datapointV_1_fu_674_p2[12]) );
  XOR2X1 U14215 ( .A(n8566), .B(n7639), .Y(datapointV_1_fu_674_p2[13]) );
  XOR2X1 U14216 ( .A(n8570), .B(n6945), .Y(datapointV_1_fu_674_p2[14]) );
  XOR2X1 U14217 ( .A(n8575), .B(n8115), .Y(datapointV_1_fu_674_p2[15]) );
  XOR2X1 U14218 ( .A(n8115), .B(n8637), .Y(datapointV_1_fu_674_p2[16]) );
  XOR2X1 U14219 ( .A(n8107), .B(n6093), .Y(datapointA_1_fu_1017_p2[1]) );
  XOR2X1 U14220 ( .A(n8554), .B(n6458), .Y(datapointA_1_fu_1017_p2[2]) );
  XOR2X1 U14221 ( .A(n8558), .B(n6946), .Y(datapointA_1_fu_1017_p2[3]) );
  XOR2X1 U14222 ( .A(n8548), .B(n7640), .Y(datapointA_1_fu_1017_p2[4]) );
  XOR2X1 U14223 ( .A(n8550), .B(n7437), .Y(datapointA_1_fu_1017_p2[5]) );
  XOR2X1 U14224 ( .A(n8553), .B(n6571), .Y(datapointA_1_fu_1017_p2[6]) );
  XOR2X1 U14225 ( .A(n8557), .B(n6164), .Y(datapointA_1_fu_1017_p2[7]) );
  XOR2X1 U14226 ( .A(n8559), .B(n6811), .Y(datapointA_1_fu_1017_p2[8]) );
  XOR2X1 U14227 ( .A(n8551), .B(n7263), .Y(datapointA_1_fu_1017_p2[9]) );
  XOR2X1 U14228 ( .A(n8555), .B(n6349), .Y(datapointA_1_fu_1017_p2[10]) );
  XOR2X1 U14229 ( .A(n8560), .B(n6686), .Y(datapointA_1_fu_1017_p2[11]) );
  XOR2X1 U14230 ( .A(n8549), .B(n7858), .Y(datapointA_1_fu_1017_p2[12]) );
  XOR2X1 U14231 ( .A(n8552), .B(n7098), .Y(datapointA_1_fu_1017_p2[13]) );
  XOR2X1 U14232 ( .A(n8556), .B(n6252), .Y(datapointA_1_fu_1017_p2[14]) );
  XOR2X1 U14233 ( .A(n8561), .B(n8408), .Y(datapointA_1_fu_1017_p2[15]) );
  XOR2X1 U14234 ( .A(n8408), .B(n8636), .Y(datapointA_1_fu_1017_p2[16]) );
  XOR2X1 U14235 ( .A(n8843), .B(p_tmp_i_reg_1556[2]), .Y(i_1_fu_620_p2[2]) );
  XOR2X1 U14236 ( .A(n8664), .B(p_tmp_i_reg_1556[3]), .Y(i_1_fu_620_p2[3]) );
  NOR3X1 U14237 ( .A(AbeatDelay_new_reg_394[16]), .B(
        AbeatDelay_new_reg_394[18]), .C(AbeatDelay_new_reg_394[17]), .Y(n11055) );
  NOR3X1 U14238 ( .A(n11048), .B(AbeatDelay_new_reg_394[20]), .C(
        AbeatDelay_new_reg_394[19]), .Y(n11054) );
  NOR3X1 U14239 ( .A(n11049), .B(AbeatDelay_new_reg_394[24]), .C(
        AbeatDelay_new_reg_394[23]), .Y(n11052) );
  NOR3X1 U14240 ( .A(n11050), .B(AbeatDelay_new_reg_394[28]), .C(
        AbeatDelay_new_reg_394[27]), .Y(n11051) );
  NAND3X1 U14241 ( .A(n11055), .B(n11054), .C(n11053), .Y(n11066) );
  AOI21X1 U14242 ( .A(n5521), .B(n11063), .C(AbeatDelay_new_reg_394[31]), .Y(
        n11065) );
  NAND3X1 U14243 ( .A(AbeatDelay_new_reg_394[6]), .B(AbeatDelay_new_reg_394[5]), .C(AbeatDelay_new_reg_394[7]), .Y(n11058) );
  NOR3X1 U14244 ( .A(AbeatDelay_new_reg_394[0]), .B(AbeatDelay_new_reg_394[2]), 
        .C(AbeatDelay_new_reg_394[1]), .Y(n11059) );
  AOI22X1 U14245 ( .A(AbeatDelay_new_reg_394[4]), .B(n10688), .C(n5754), .D(
        AbeatDelay_new_reg_394[3]), .Y(n11061) );
  NAND3X1 U14246 ( .A(n11063), .B(n8308), .C(n5757), .Y(n11064) );
  AOI22X1 U14247 ( .A(n5562), .B(n10741), .C(n5737), .D(n5755), .Y(n11067) );
  NOR3X1 U14248 ( .A(AbeatDelay_new_reg_394[16]), .B(
        AbeatDelay_new_reg_394[18]), .C(AbeatDelay_new_reg_394[17]), .Y(n11075) );
  NOR3X1 U14249 ( .A(n11068), .B(AbeatDelay_new_reg_394[20]), .C(
        AbeatDelay_new_reg_394[19]), .Y(n11074) );
  NOR3X1 U14250 ( .A(n11069), .B(AbeatDelay_new_reg_394[24]), .C(
        AbeatDelay_new_reg_394[23]), .Y(n11072) );
  NOR3X1 U14251 ( .A(n11070), .B(AbeatDelay_new_reg_394[28]), .C(
        AbeatDelay_new_reg_394[27]), .Y(n11071) );
  NAND3X1 U14252 ( .A(n11075), .B(n11074), .C(n11073), .Y(n11084) );
  AOI21X1 U14253 ( .A(AbeatDelay_new_reg_394[9]), .B(AbeatDelay_new_reg_394[8]), .C(n11062), .Y(n11076) );
  AOI21X1 U14254 ( .A(n5521), .B(n11081), .C(AbeatDelay_new_reg_394[31]), .Y(
        n11083) );
  NOR3X1 U14255 ( .A(AbeatDelay_new_reg_394[0]), .B(AbeatDelay_new_reg_394[3]), 
        .C(AbeatDelay_new_reg_394[1]), .Y(n11077) );
  OAI21X1 U14256 ( .A(AbeatDelay_new_reg_394[2]), .B(AbeatDelay_new_reg_394[3]), .C(n10676), .Y(n11078) );
  NOR3X1 U14257 ( .A(AbeatDelay_new_reg_394[4]), .B(AbeatDelay_new_reg_394[6]), 
        .C(AbeatDelay_new_reg_394[5]), .Y(n11079) );
  AOI22X1 U14258 ( .A(n10675), .B(AbeatDelay_new_reg_394[7]), .C(
        AbeatDelay_new_reg_394[7]), .D(n10685), .Y(n11080) );
  NAND3X1 U14259 ( .A(n11081), .B(n8308), .C(n5758), .Y(n11082) );
  AOI22X1 U14260 ( .A(n5563), .B(n10741), .C(n5738), .D(n5756), .Y(n11085) );
  OAI21X1 U14261 ( .A(VbeatDelay_new_1_reg_326[14]), .B(n10707), .C(n8074), 
        .Y(n11086) );
  NAND3X1 U14262 ( .A(n11097), .B(n11087), .C(n10487), .Y(n11105) );
  OAI21X1 U14263 ( .A(VbeatDelay_new_1_reg_326[10]), .B(n10699), .C(n8075), 
        .Y(n11088) );
  NAND3X1 U14264 ( .A(n8075), .B(n10699), .C(VbeatDelay_new_1_reg_326[10]), 
        .Y(n11090) );
  OAI21X1 U14265 ( .A(AbeatDelay_new_reg_394[11]), .B(n10480), .C(n7208), .Y(
        n11094) );
  NOR3X1 U14266 ( .A(n8089), .B(AbeatDelay_new_reg_394[8]), .C(n10472), .Y(
        n11091) );
  NAND3X1 U14267 ( .A(n10471), .B(n7592), .C(n10477), .Y(n11093) );
  OAI21X1 U14268 ( .A(n10476), .B(n11094), .C(n7591), .Y(n11103) );
  NAND3X1 U14269 ( .A(n8074), .B(n10707), .C(VbeatDelay_new_1_reg_326[14]), 
        .Y(n11096) );
  OAI21X1 U14270 ( .A(AbeatDelay_new_reg_394[15]), .B(n10491), .C(n4820), .Y(
        n11101) );
  NAND3X1 U14271 ( .A(n11097), .B(n10703), .C(VbeatDelay_new_1_reg_326[12]), 
        .Y(n11099) );
  NAND3X1 U14272 ( .A(n5452), .B(n8002), .C(n10488), .Y(n11100) );
  OAI21X1 U14273 ( .A(n10487), .B(n11101), .C(n4821), .Y(n11102) );
  OAI21X1 U14274 ( .A(n8307), .B(n11103), .C(n11102), .Y(n11104) );
  AOI21X1 U14275 ( .A(AbeatDelay_new_reg_394[8]), .B(n10472), .C(n8089), .Y(
        n11107) );
  NAND3X1 U14276 ( .A(n10476), .B(n10482), .C(n5861), .Y(n11126) );
  AOI21X1 U14277 ( .A(AbeatDelay_new_reg_394[1]), .B(n10454), .C(
        AbeatDelay_new_reg_394[0]), .Y(n11108) );
  AOI22X1 U14278 ( .A(VbeatDelay_new_1_reg_326[1]), .B(n10679), .C(n8013), .D(
        VbeatDelay_new_1_reg_326[0]), .Y(n11111) );
  NAND3X1 U14279 ( .A(n8083), .B(n10681), .C(VbeatDelay_new_1_reg_326[2]), .Y(
        n11109) );
  OAI21X1 U14280 ( .A(AbeatDelay_new_reg_394[3]), .B(n10459), .C(n4822), .Y(
        n11110) );
  OAI21X1 U14281 ( .A(VbeatDelay_new_1_reg_326[6]), .B(n10691), .C(n8084), .Y(
        n11121) );
  AOI21X1 U14282 ( .A(n8012), .B(n10456), .C(n11121), .Y(n11124) );
  OAI21X1 U14283 ( .A(VbeatDelay_new_1_reg_326[2]), .B(n10681), .C(n8083), .Y(
        n11114) );
  OAI21X1 U14284 ( .A(VbeatDelay_new_1_reg_326[4]), .B(n10686), .C(n11118), 
        .Y(n11113) );
  AOI21X1 U14285 ( .A(n10456), .B(n11114), .C(n11113), .Y(n11123) );
  NAND3X1 U14286 ( .A(n8084), .B(n10691), .C(VbeatDelay_new_1_reg_326[6]), .Y(
        n11116) );
  OAI21X1 U14287 ( .A(AbeatDelay_new_reg_394[7]), .B(n10468), .C(n4823), .Y(
        n11117) );
  AOI22X1 U14288 ( .A(VbeatDelay_new_1_reg_326[5]), .B(n10689), .C(n11119), 
        .D(VbeatDelay_new_1_reg_326[4]), .Y(n11120) );
  AOI22X1 U14289 ( .A(n10465), .B(n11121), .C(n8247), .D(n10465), .Y(n11122)
         );
  AOI21X1 U14290 ( .A(n5522), .B(n5501), .C(n5295), .Y(n11125) );
  AOI22X1 U14291 ( .A(n10470), .B(n5551), .C(n5739), .D(n10470), .Y(n11127) );
  NAND3X1 U14292 ( .A(n11155), .B(n11128), .C(n5759), .Y(n11174) );
  OAI21X1 U14293 ( .A(VbeatDelay_new_1_reg_326[18]), .B(n10715), .C(n8080), 
        .Y(n11158) );
  OAI21X1 U14294 ( .A(VbeatDelay_new_1_reg_326[22]), .B(n10723), .C(n8079), 
        .Y(n11165) );
  NAND3X1 U14295 ( .A(n11162), .B(n11129), .C(n10508), .Y(n11130) );
  OAI21X1 U14296 ( .A(VbeatDelay_new_1_reg_326[26]), .B(n10731), .C(n8073), 
        .Y(n11134) );
  OAI21X1 U14297 ( .A(VbeatDelay_new_1_reg_326[30]), .B(n10739), .C(n8325), 
        .Y(n11131) );
  NAND3X1 U14298 ( .A(n11144), .B(n11132), .C(n10529), .Y(n11151) );
  OAI21X1 U14299 ( .A(n10727), .B(VbeatDelay_new_1_reg_326[24]), .C(n11137), 
        .Y(n11133) );
  NOR3X1 U14300 ( .A(n11134), .B(n8099), .C(n11133), .Y(n11171) );
  NAND3X1 U14301 ( .A(n10497), .B(n10503), .C(n11171), .Y(n11173) );
  NAND3X1 U14302 ( .A(n8073), .B(n10731), .C(VbeatDelay_new_1_reg_326[26]), 
        .Y(n11136) );
  OAI21X1 U14303 ( .A(AbeatDelay_new_reg_394[27]), .B(n10523), .C(n4824), .Y(
        n11141) );
  NAND3X1 U14304 ( .A(n11137), .B(n10727), .C(VbeatDelay_new_1_reg_326[24]), 
        .Y(n11139) );
  NAND3X1 U14305 ( .A(n5453), .B(n5571), .C(n10520), .Y(n11140) );
  OAI21X1 U14306 ( .A(n10519), .B(n11141), .C(n4825), .Y(n11150) );
  NAND3X1 U14307 ( .A(n8325), .B(n10739), .C(VbeatDelay_new_1_reg_326[30]), 
        .Y(n11143) );
  OAI21X1 U14308 ( .A(VbeatDelay_new_1_reg_326[31]), .B(n10741), .C(n4826), 
        .Y(n11148) );
  NAND3X1 U14309 ( .A(n11144), .B(n10735), .C(VbeatDelay_new_1_reg_326[28]), 
        .Y(n11146) );
  NAND3X1 U14310 ( .A(n5454), .B(n7789), .C(n10530), .Y(n11147) );
  OAI21X1 U14311 ( .A(n10529), .B(n11148), .C(n4827), .Y(n11149) );
  OAI21X1 U14312 ( .A(n8099), .B(n11150), .C(n11149), .Y(n11170) );
  NAND3X1 U14313 ( .A(n8080), .B(n10715), .C(VbeatDelay_new_1_reg_326[18]), 
        .Y(n11153) );
  OAI21X1 U14314 ( .A(AbeatDelay_new_reg_394[19]), .B(n10501), .C(n4828), .Y(
        n11154) );
  AOI22X1 U14315 ( .A(VbeatDelay_new_1_reg_326[17]), .B(n10713), .C(n11156), 
        .D(VbeatDelay_new_1_reg_326[16]), .Y(n11157) );
  AOI22X1 U14316 ( .A(n10498), .B(n11158), .C(n7596), .D(n10498), .Y(n11167)
         );
  NAND3X1 U14317 ( .A(n8079), .B(n10723), .C(VbeatDelay_new_1_reg_326[22]), 
        .Y(n11160) );
  OAI21X1 U14318 ( .A(AbeatDelay_new_reg_394[23]), .B(n10512), .C(n4829), .Y(
        n11161) );
  AOI22X1 U14319 ( .A(VbeatDelay_new_1_reg_326[21]), .B(n10721), .C(n11163), 
        .D(VbeatDelay_new_1_reg_326[20]), .Y(n11164) );
  AOI22X1 U14320 ( .A(n10509), .B(n11165), .C(n7407), .D(n10509), .Y(n11166)
         );
  AOI21X1 U14321 ( .A(n7595), .B(n10503), .C(n7406), .Y(n11168) );
  OAI21X1 U14322 ( .A(n11171), .B(n11170), .C(n4927), .Y(n11172) );
  OAI21X1 U14323 ( .A(n5533), .B(n5700), .C(n11172), .Y(N503) );
  XOR2X1 U14324 ( .A(\add_1121/carry[31] ), .B(recentABools_len[31]), .Y(
        CircularBuffer_len_read_assign_2_fu_1085_p2[31]) );
  XOR2X1 U14325 ( .A(\add_1125/carry[31] ), .B(recentVBools_len[31]), .Y(
        CircularBuffer_len_read_assign_fu_772_p2[31]) );
  OAI21X1 U14326 ( .A(n11204), .B(n7860), .C(n5910), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[10]) );
  OAI21X1 U14327 ( .A(n11175), .B(n8399), .C(n7827), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[11]) );
  OAI21X1 U14328 ( .A(n11176), .B(n7439), .C(n5911), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[12]) );
  OAI21X1 U14329 ( .A(n11177), .B(n7642), .C(n5912), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[13]) );
  OAI21X1 U14330 ( .A(n11178), .B(n8103), .C(n7831), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[14]) );
  OAI21X1 U14331 ( .A(n11179), .B(n8114), .C(n7621), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[15]) );
  OAI21X1 U14332 ( .A(n11180), .B(n6254), .C(n5913), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[16]) );
  OAI21X1 U14333 ( .A(n11181), .B(n6351), .C(n5914), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[17]) );
  OAI21X1 U14334 ( .A(n11182), .B(n7443), .C(n5915), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[18]) );
  OAI21X1 U14335 ( .A(n11183), .B(n7864), .C(n5916), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[19]) );
  OAI21X1 U14336 ( .A(n8392), .B(n10539), .C(n8055), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[1]) );
  OAI21X1 U14337 ( .A(n11185), .B(n6460), .C(n5917), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[20]) );
  OAI21X1 U14338 ( .A(n11186), .B(n7265), .C(n5918), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[21]) );
  OAI21X1 U14339 ( .A(n11187), .B(n7100), .C(n5919), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[22]) );
  OAI21X1 U14340 ( .A(n11188), .B(n8401), .C(n7829), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[23]) );
  OAI21X1 U14341 ( .A(n11189), .B(n6573), .C(n5920), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[24]) );
  OAI21X1 U14342 ( .A(n11190), .B(n6948), .C(n5921), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[25]) );
  OAI21X1 U14343 ( .A(n11191), .B(n6813), .C(n5922), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[26]) );
  OAI21X1 U14344 ( .A(n11192), .B(n7646), .C(n5923), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[27]) );
  OAI21X1 U14345 ( .A(n11193), .B(n6688), .C(n5924), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[28]) );
  OAI21X1 U14346 ( .A(n11194), .B(n6166), .C(n8386), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[29]) );
  OAI21X1 U14347 ( .A(n11184), .B(n10538), .C(n8298), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[2]) );
  XNOR2X1 U14348 ( .A(n2238), .B(n8386), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[30]) );
  XNOR2X1 U14349 ( .A(n2401), .B(n11197), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[31]) );
  OAI21X1 U14350 ( .A(n11195), .B(n10537), .C(n8053), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[3]) );
  OAI21X1 U14351 ( .A(n11198), .B(n10536), .C(n8296), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[4]) );
  OAI21X1 U14352 ( .A(n11199), .B(n7441), .C(n5908), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[5]) );
  OAI21X1 U14353 ( .A(n11200), .B(n7644), .C(n5909), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[6]) );
  OAI21X1 U14354 ( .A(n11201), .B(n8112), .C(n7619), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[7]) );
  OAI21X1 U14355 ( .A(n11202), .B(n8407), .C(n8051), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[8]) );
  OAI21X1 U14356 ( .A(n11203), .B(n7862), .C(n7617), .Y(
        CircularBuffer_len_write_assig_2_fu_1142_p2[9]) );
  OAI21X1 U14357 ( .A(n11234), .B(n7859), .C(n5927), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[10]) );
  OAI21X1 U14358 ( .A(n11205), .B(n8398), .C(n7826), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[11]) );
  OAI21X1 U14359 ( .A(n11206), .B(n7438), .C(n5928), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[12]) );
  OAI21X1 U14360 ( .A(n11207), .B(n7641), .C(n5929), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[13]) );
  OAI21X1 U14361 ( .A(n11208), .B(n8102), .C(n7830), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[14]) );
  OAI21X1 U14362 ( .A(n11209), .B(n8113), .C(n7620), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[15]) );
  OAI21X1 U14363 ( .A(n11210), .B(n6253), .C(n5930), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[16]) );
  OAI21X1 U14364 ( .A(n11211), .B(n6350), .C(n5931), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[17]) );
  OAI21X1 U14365 ( .A(n11212), .B(n7442), .C(n5932), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[18]) );
  OAI21X1 U14366 ( .A(n11213), .B(n7863), .C(n5933), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[19]) );
  OAI21X1 U14367 ( .A(n8391), .B(n10074), .C(n8054), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[1]) );
  OAI21X1 U14368 ( .A(n11215), .B(n6459), .C(n5934), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[20]) );
  OAI21X1 U14369 ( .A(n11216), .B(n7264), .C(n5935), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[21]) );
  OAI21X1 U14370 ( .A(n11217), .B(n7099), .C(n5936), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[22]) );
  OAI21X1 U14371 ( .A(n11218), .B(n8400), .C(n7828), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[23]) );
  OAI21X1 U14372 ( .A(n11219), .B(n6572), .C(n5937), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[24]) );
  OAI21X1 U14373 ( .A(n11220), .B(n6947), .C(n5938), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[25]) );
  OAI21X1 U14374 ( .A(n11221), .B(n6812), .C(n5939), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[26]) );
  OAI21X1 U14375 ( .A(n11222), .B(n7645), .C(n5940), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[27]) );
  OAI21X1 U14376 ( .A(n11223), .B(n6687), .C(n5941), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[28]) );
  OAI21X1 U14377 ( .A(n11224), .B(n6165), .C(n8385), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[29]) );
  OAI21X1 U14378 ( .A(n11214), .B(n10073), .C(n8297), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[2]) );
  XNOR2X1 U14379 ( .A(n2734), .B(n8385), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[30]) );
  XNOR2X1 U14380 ( .A(n2862), .B(n11227), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[31]) );
  OAI21X1 U14381 ( .A(n11225), .B(n10072), .C(n8052), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[3]) );
  OAI21X1 U14382 ( .A(n11228), .B(n10071), .C(n8295), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[4]) );
  OAI21X1 U14383 ( .A(n11229), .B(n7440), .C(n5925), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[5]) );
  OAI21X1 U14384 ( .A(n11230), .B(n7643), .C(n5926), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[6]) );
  OAI21X1 U14385 ( .A(n11231), .B(n8111), .C(n7618), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[7]) );
  OAI21X1 U14386 ( .A(n11232), .B(n8406), .C(n8050), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[8]) );
  OAI21X1 U14387 ( .A(n11233), .B(n7861), .C(n7616), .Y(
        CircularBuffer_len_write_assig_fu_817_p2[9]) );
  OAI21X1 U14388 ( .A(n9900), .B(n9899), .C(n8299), .Y(i_fu_607_p2[1]) );
  OAI21X1 U14389 ( .A(n11235), .B(n9898), .C(n8056), .Y(i_fu_607_p2[2]) );
  NOR3X1 U14390 ( .A(p_tmp_i_reg_1556[23]), .B(p_tmp_i_reg_1556[25]), .C(
        p_tmp_i_reg_1556[24]), .Y(n11242) );
  NOR3X1 U14391 ( .A(n11236), .B(p_tmp_i_reg_1556[27]), .C(
        p_tmp_i_reg_1556[26]), .Y(n11241) );
  NOR3X1 U14392 ( .A(p_tmp_i_reg_1556[30]), .B(p_tmp_i_reg_1556[5]), .C(
        p_tmp_i_reg_1556[4]), .Y(n11239) );
  NOR3X1 U14393 ( .A(n11237), .B(p_tmp_i_reg_1556[7]), .C(p_tmp_i_reg_1556[6]), 
        .Y(n11238) );
  NAND3X1 U14394 ( .A(n11242), .B(n11241), .C(n11240), .Y(n11252) );
  NOR3X1 U14395 ( .A(p_tmp_i_reg_1556[16]), .B(p_tmp_i_reg_1556[18]), .C(
        p_tmp_i_reg_1556[17]), .Y(n11243) );
  NAND3X1 U14396 ( .A(n7590), .B(n8240), .C(n11243), .Y(n11251) );
  NOR3X1 U14397 ( .A(n11247), .B(p_tmp_i_reg_1556[13]), .C(
        p_tmp_i_reg_1556[12]), .Y(n11248) );
  NAND3X1 U14398 ( .A(n8048), .B(n11254), .C(n11248), .Y(n11250) );
  NOR3X1 U14399 ( .A(n7804), .B(n7805), .C(n8047), .Y(n11253) );
  XOR2X1 U14400 ( .A(p_tmp_i_reg_1556[31]), .B(n11253), .Y(i_fu_607_p2_31) );
  OAI21X1 U14401 ( .A(n11246), .B(n9897), .C(n8384), .Y(i_fu_607_p2[3]) );
  XNOR2X1 U14402 ( .A(p_tmp_i_reg_1556[4]), .B(n8384), .Y(i_fu_607_p2[4]) );
  OAI21X1 U14403 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[5]), .B(n10639), .C(\sub_1255/carry[5] ), .Y(n11255) );
  AOI21X1 U14404 ( .A(n10639), .B(CircularBuffer_head_i_read_ass_1_reg_1719[5]), .C(n10304), .Y(n11257) );
  AOI21X1 U14405 ( .A(n10333), .B(n8370), .C(
        CircularBuffer_len_write_assig_2_reg_1729[6]), .Y(n11256) );
  OAI21X1 U14406 ( .A(n8370), .B(n10333), .C(n10303), .Y(n11258) );
  OAI21X1 U14407 ( .A(CircularBuffer_len_write_assig_2_reg_1729[7]), .B(n8008), 
        .C(n8009), .Y(n11262) );
  AOI21X1 U14408 ( .A(n10334), .B(n10302), .C(
        CircularBuffer_len_write_assig_2_reg_1729[8]), .Y(n11261) );
  AOI21X1 U14409 ( .A(n11262), .B(CircularBuffer_head_i_read_ass_1_reg_1719[8]), .C(n5309), .Y(n11264) );
  AOI21X1 U14410 ( .A(n10335), .B(n7854), .C(
        CircularBuffer_len_write_assig_2_reg_1729[9]), .Y(n11263) );
  OAI21X1 U14411 ( .A(n7854), .B(n10335), .C(n10301), .Y(n11266) );
  AOI21X1 U14412 ( .A(n10336), .B(n10300), .C(
        CircularBuffer_len_write_assig_2_reg_1729[10]), .Y(n11265) );
  AOI21X1 U14413 ( .A(n11266), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[10]), .C(n5310), .Y(n11268)
         );
  AOI21X1 U14414 ( .A(n10337), .B(n5975), .C(
        CircularBuffer_len_write_assig_2_reg_1729[11]), .Y(n11267) );
  OAI21X1 U14415 ( .A(n5975), .B(n10337), .C(n10299), .Y(n11270) );
  AOI21X1 U14416 ( .A(n10338), .B(n10298), .C(
        CircularBuffer_len_write_assig_2_reg_1729[12]), .Y(n11269) );
  AOI21X1 U14417 ( .A(n11270), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[12]), .C(n5311), .Y(n11272)
         );
  AOI21X1 U14418 ( .A(n10339), .B(n5976), .C(
        CircularBuffer_len_write_assig_2_reg_1729[13]), .Y(n11271) );
  OAI21X1 U14419 ( .A(n5976), .B(n10339), .C(n10297), .Y(n11274) );
  AOI21X1 U14420 ( .A(n10340), .B(n10296), .C(
        CircularBuffer_len_write_assig_2_reg_1729[14]), .Y(n11273) );
  AOI21X1 U14421 ( .A(n11274), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[14]), .C(n5312), .Y(n11276)
         );
  AOI21X1 U14422 ( .A(n10341), .B(n5977), .C(
        CircularBuffer_len_write_assig_2_reg_1729[15]), .Y(n11275) );
  OAI21X1 U14423 ( .A(n5977), .B(n10341), .C(n10295), .Y(n11278) );
  AOI21X1 U14424 ( .A(n10342), .B(n10294), .C(
        CircularBuffer_len_write_assig_2_reg_1729[16]), .Y(n11277) );
  AOI21X1 U14425 ( .A(n11278), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[16]), .C(n5313), .Y(n11280)
         );
  AOI21X1 U14426 ( .A(n10343), .B(n5978), .C(
        CircularBuffer_len_write_assig_2_reg_1729[17]), .Y(n11279) );
  OAI21X1 U14427 ( .A(n5978), .B(n10343), .C(n10293), .Y(n11282) );
  AOI21X1 U14428 ( .A(n10344), .B(n10292), .C(
        CircularBuffer_len_write_assig_2_reg_1729[18]), .Y(n11281) );
  AOI21X1 U14429 ( .A(n11282), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[18]), .C(n5314), .Y(n11284)
         );
  AOI21X1 U14430 ( .A(n10345), .B(n5979), .C(
        CircularBuffer_len_write_assig_2_reg_1729[19]), .Y(n11283) );
  OAI21X1 U14431 ( .A(n5979), .B(n10345), .C(n10291), .Y(n11286) );
  AOI21X1 U14432 ( .A(n10346), .B(n10290), .C(
        CircularBuffer_len_write_assig_2_reg_1729[20]), .Y(n11285) );
  AOI21X1 U14433 ( .A(n11286), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[20]), .C(n5315), .Y(n11288)
         );
  AOI21X1 U14434 ( .A(n10347), .B(n5980), .C(
        CircularBuffer_len_write_assig_2_reg_1729[21]), .Y(n11287) );
  OAI21X1 U14435 ( .A(n5980), .B(n10347), .C(n10289), .Y(n11290) );
  AOI21X1 U14436 ( .A(n10348), .B(n10288), .C(
        CircularBuffer_len_write_assig_2_reg_1729[22]), .Y(n11289) );
  AOI21X1 U14437 ( .A(n11290), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[22]), .C(n5316), .Y(n11292)
         );
  AOI21X1 U14438 ( .A(n10349), .B(n5981), .C(
        CircularBuffer_len_write_assig_2_reg_1729[23]), .Y(n11291) );
  OAI21X1 U14439 ( .A(n5981), .B(n10349), .C(n10287), .Y(n11294) );
  AOI21X1 U14440 ( .A(n10350), .B(n10286), .C(
        CircularBuffer_len_write_assig_2_reg_1729[24]), .Y(n11293) );
  AOI21X1 U14441 ( .A(n11294), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[24]), .C(n5317), .Y(n11296)
         );
  AOI21X1 U14442 ( .A(n10351), .B(n5982), .C(
        CircularBuffer_len_write_assig_2_reg_1729[25]), .Y(n11295) );
  OAI21X1 U14443 ( .A(n5982), .B(n10351), .C(n10285), .Y(n11298) );
  AOI21X1 U14444 ( .A(n10352), .B(n10284), .C(
        CircularBuffer_len_write_assig_2_reg_1729[26]), .Y(n11297) );
  AOI21X1 U14445 ( .A(n11298), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[26]), .C(n5318), .Y(n11300)
         );
  AOI21X1 U14446 ( .A(n10353), .B(n5983), .C(
        CircularBuffer_len_write_assig_2_reg_1729[27]), .Y(n11299) );
  OAI21X1 U14447 ( .A(n5983), .B(n10353), .C(n10283), .Y(n11302) );
  AOI21X1 U14448 ( .A(n10354), .B(n10282), .C(
        CircularBuffer_len_write_assig_2_reg_1729[28]), .Y(n11301) );
  AOI21X1 U14449 ( .A(n11302), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[28]), .C(n5319), .Y(n11303)
         );
  AOI21X1 U14450 ( .A(n10355), .B(n8098), .C(
        CircularBuffer_len_write_assig_2_reg_1729[29]), .Y(n11304) );
  AOI21X1 U14451 ( .A(n10281), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[29]), .C(n8097), .Y(n11306)
         );
  AOI21X1 U14452 ( .A(n10356), .B(n8096), .C(
        CircularBuffer_len_write_assig_2_reg_1729[30]), .Y(n11305) );
  OAI21X1 U14453 ( .A(n8096), .B(n10356), .C(n10280), .Y(\sub_1255/carry[31] )
         );
  OAI21X1 U14454 ( .A(CircularBuffer_head_i_read_ass_reg_1624[5]), .B(n10083), 
        .C(\sub_1263/carry[5] ), .Y(n11307) );
  AOI21X1 U14455 ( .A(n10083), .B(CircularBuffer_head_i_read_ass_reg_1624[5]), 
        .C(n9990), .Y(n11309) );
  AOI21X1 U14456 ( .A(n10026), .B(n8369), .C(
        CircularBuffer_len_read_assign_1_reg_1616[6]), .Y(n11308) );
  OAI21X1 U14457 ( .A(n8369), .B(n10026), .C(n9989), .Y(n11310) );
  OAI21X1 U14458 ( .A(CircularBuffer_len_read_assign_1_reg_1616[7]), .B(n8006), 
        .C(n8007), .Y(n11314) );
  AOI21X1 U14459 ( .A(n10027), .B(n9988), .C(
        CircularBuffer_len_read_assign_1_reg_1616[8]), .Y(n11313) );
  AOI21X1 U14460 ( .A(n11314), .B(CircularBuffer_head_i_read_ass_reg_1624[8]), 
        .C(n5320), .Y(n11316) );
  AOI21X1 U14461 ( .A(n10028), .B(n7852), .C(
        CircularBuffer_len_read_assign_1_reg_1616[9]), .Y(n11315) );
  OAI21X1 U14462 ( .A(n7852), .B(n10028), .C(n9987), .Y(n11318) );
  AOI21X1 U14463 ( .A(n10029), .B(n9986), .C(
        CircularBuffer_len_read_assign_1_reg_1616[10]), .Y(n11317) );
  AOI21X1 U14464 ( .A(n11318), .B(CircularBuffer_head_i_read_ass_reg_1624[10]), 
        .C(n5321), .Y(n11320) );
  AOI21X1 U14465 ( .A(n10030), .B(n5984), .C(
        CircularBuffer_len_read_assign_1_reg_1616[11]), .Y(n11319) );
  OAI21X1 U14466 ( .A(n5984), .B(n10030), .C(n9985), .Y(n11322) );
  AOI21X1 U14467 ( .A(n10031), .B(n9984), .C(
        CircularBuffer_len_read_assign_1_reg_1616[12]), .Y(n11321) );
  AOI21X1 U14468 ( .A(n11322), .B(CircularBuffer_head_i_read_ass_reg_1624[12]), 
        .C(n5322), .Y(n11324) );
  AOI21X1 U14469 ( .A(n10032), .B(n5985), .C(
        CircularBuffer_len_read_assign_1_reg_1616[13]), .Y(n11323) );
  OAI21X1 U14470 ( .A(n5985), .B(n10032), .C(n9983), .Y(n11326) );
  AOI21X1 U14471 ( .A(n10033), .B(n9982), .C(
        CircularBuffer_len_read_assign_1_reg_1616[14]), .Y(n11325) );
  AOI21X1 U14472 ( .A(n11326), .B(CircularBuffer_head_i_read_ass_reg_1624[14]), 
        .C(n5323), .Y(n11328) );
  AOI21X1 U14473 ( .A(n10034), .B(n5986), .C(
        CircularBuffer_len_read_assign_1_reg_1616[15]), .Y(n11327) );
  OAI21X1 U14474 ( .A(n5986), .B(n10034), .C(n9981), .Y(n11330) );
  AOI21X1 U14475 ( .A(n10035), .B(n9980), .C(
        CircularBuffer_len_read_assign_1_reg_1616[16]), .Y(n11329) );
  AOI21X1 U14476 ( .A(n11330), .B(CircularBuffer_head_i_read_ass_reg_1624[16]), 
        .C(n5324), .Y(n11332) );
  AOI21X1 U14477 ( .A(n10036), .B(n5987), .C(
        CircularBuffer_len_read_assign_1_reg_1616[17]), .Y(n11331) );
  OAI21X1 U14478 ( .A(n5987), .B(n10036), .C(n9979), .Y(n11334) );
  AOI21X1 U14479 ( .A(n10037), .B(n9978), .C(
        CircularBuffer_len_read_assign_1_reg_1616[18]), .Y(n11333) );
  AOI21X1 U14480 ( .A(n11334), .B(CircularBuffer_head_i_read_ass_reg_1624[18]), 
        .C(n5325), .Y(n11336) );
  AOI21X1 U14481 ( .A(n10038), .B(n5988), .C(
        CircularBuffer_len_read_assign_1_reg_1616[19]), .Y(n11335) );
  OAI21X1 U14482 ( .A(n5988), .B(n10038), .C(n9977), .Y(n11338) );
  AOI21X1 U14483 ( .A(n10039), .B(n9976), .C(
        CircularBuffer_len_read_assign_1_reg_1616[20]), .Y(n11337) );
  AOI21X1 U14484 ( .A(n11338), .B(CircularBuffer_head_i_read_ass_reg_1624[20]), 
        .C(n5326), .Y(n11340) );
  AOI21X1 U14485 ( .A(n10040), .B(n5989), .C(
        CircularBuffer_len_read_assign_1_reg_1616[21]), .Y(n11339) );
  OAI21X1 U14486 ( .A(n5989), .B(n10040), .C(n9975), .Y(n11342) );
  AOI21X1 U14487 ( .A(n10041), .B(n9974), .C(
        CircularBuffer_len_read_assign_1_reg_1616[22]), .Y(n11341) );
  AOI21X1 U14488 ( .A(n11342), .B(CircularBuffer_head_i_read_ass_reg_1624[22]), 
        .C(n5327), .Y(n11344) );
  AOI21X1 U14489 ( .A(n10042), .B(n5990), .C(
        CircularBuffer_len_read_assign_1_reg_1616[23]), .Y(n11343) );
  OAI21X1 U14490 ( .A(n5990), .B(n10042), .C(n9973), .Y(n11346) );
  AOI21X1 U14491 ( .A(n10043), .B(n9972), .C(
        CircularBuffer_len_read_assign_1_reg_1616[24]), .Y(n11345) );
  AOI21X1 U14492 ( .A(n11346), .B(CircularBuffer_head_i_read_ass_reg_1624[24]), 
        .C(n5328), .Y(n11348) );
  AOI21X1 U14493 ( .A(n10044), .B(n5991), .C(
        CircularBuffer_len_read_assign_1_reg_1616[25]), .Y(n11347) );
  OAI21X1 U14494 ( .A(n5991), .B(n10044), .C(n9971), .Y(n11350) );
  AOI21X1 U14495 ( .A(n10045), .B(n9970), .C(
        CircularBuffer_len_read_assign_1_reg_1616[26]), .Y(n11349) );
  AOI21X1 U14496 ( .A(n11350), .B(CircularBuffer_head_i_read_ass_reg_1624[26]), 
        .C(n5329), .Y(n11352) );
  AOI21X1 U14497 ( .A(n10046), .B(n8092), .C(
        CircularBuffer_len_read_assign_1_reg_1616[27]), .Y(n11351) );
  OAI21X1 U14498 ( .A(n8092), .B(n10046), .C(n9969), .Y(n11354) );
  AOI21X1 U14499 ( .A(n10047), .B(n9968), .C(
        CircularBuffer_len_read_assign_1_reg_1616[28]), .Y(n11353) );
  AOI21X1 U14500 ( .A(n11354), .B(CircularBuffer_head_i_read_ass_reg_1624[28]), 
        .C(n5330), .Y(n11355) );
  AOI21X1 U14501 ( .A(n10048), .B(n8365), .C(
        CircularBuffer_len_read_assign_1_reg_1616[29]), .Y(n11356) );
  AOI21X1 U14502 ( .A(n9967), .B(CircularBuffer_head_i_read_ass_reg_1624[29]), 
        .C(n8364), .Y(n11358) );
  AOI21X1 U14503 ( .A(n10049), .B(n8363), .C(
        CircularBuffer_len_read_assign_1_reg_1616[30]), .Y(n11357) );
  OAI21X1 U14504 ( .A(n8363), .B(n10049), .C(n9966), .Y(\sub_1263/carry[31] )
         );
  OAI21X1 U14505 ( .A(CircularBuffer_head_i_read_ass_reg_1624[5]), .B(n10144), 
        .C(\sub_1269/carry[5] ), .Y(n11359) );
  AOI21X1 U14506 ( .A(n10144), .B(CircularBuffer_head_i_read_ass_reg_1624[5]), 
        .C(n10022), .Y(n11361) );
  AOI21X1 U14507 ( .A(n10026), .B(n8090), .C(
        CircularBuffer_len_write_assig_reg_1634[6]), .Y(n11360) );
  OAI21X1 U14508 ( .A(n8090), .B(n10026), .C(n10021), .Y(n11362) );
  OAI21X1 U14509 ( .A(CircularBuffer_len_write_assig_reg_1634[7]), .B(n8241), 
        .C(n8242), .Y(n11366) );
  AOI21X1 U14510 ( .A(n10027), .B(n10020), .C(
        CircularBuffer_len_write_assig_reg_1634[8]), .Y(n11365) );
  AOI21X1 U14511 ( .A(n11366), .B(CircularBuffer_head_i_read_ass_reg_1624[8]), 
        .C(n5331), .Y(n11368) );
  AOI21X1 U14512 ( .A(n10028), .B(n7635), .C(
        CircularBuffer_len_write_assig_reg_1634[9]), .Y(n11367) );
  OAI21X1 U14513 ( .A(n7635), .B(n10028), .C(n10019), .Y(n11370) );
  AOI21X1 U14514 ( .A(n10029), .B(n10018), .C(
        CircularBuffer_len_write_assig_reg_1634[10]), .Y(n11369) );
  AOI21X1 U14515 ( .A(n11370), .B(CircularBuffer_head_i_read_ass_reg_1624[10]), 
        .C(n5332), .Y(n11372) );
  AOI21X1 U14516 ( .A(n10030), .B(n5992), .C(
        CircularBuffer_len_write_assig_reg_1634[11]), .Y(n11371) );
  OAI21X1 U14517 ( .A(n5992), .B(n10030), .C(n10017), .Y(n11374) );
  AOI21X1 U14518 ( .A(n10031), .B(n10016), .C(
        CircularBuffer_len_write_assig_reg_1634[12]), .Y(n11373) );
  AOI21X1 U14519 ( .A(n11374), .B(CircularBuffer_head_i_read_ass_reg_1624[12]), 
        .C(n5333), .Y(n11376) );
  AOI21X1 U14520 ( .A(n10032), .B(n5993), .C(
        CircularBuffer_len_write_assig_reg_1634[13]), .Y(n11375) );
  OAI21X1 U14521 ( .A(n5993), .B(n10032), .C(n10015), .Y(n11378) );
  AOI21X1 U14522 ( .A(n10033), .B(n10014), .C(
        CircularBuffer_len_write_assig_reg_1634[14]), .Y(n11377) );
  AOI21X1 U14523 ( .A(n11378), .B(CircularBuffer_head_i_read_ass_reg_1624[14]), 
        .C(n5334), .Y(n11380) );
  AOI21X1 U14524 ( .A(n10034), .B(n5994), .C(
        CircularBuffer_len_write_assig_reg_1634[15]), .Y(n11379) );
  OAI21X1 U14525 ( .A(n5994), .B(n10034), .C(n10013), .Y(n11382) );
  AOI21X1 U14526 ( .A(n10035), .B(n10012), .C(
        CircularBuffer_len_write_assig_reg_1634[16]), .Y(n11381) );
  AOI21X1 U14527 ( .A(n11382), .B(CircularBuffer_head_i_read_ass_reg_1624[16]), 
        .C(n5335), .Y(n11384) );
  AOI21X1 U14528 ( .A(n10036), .B(n5995), .C(
        CircularBuffer_len_write_assig_reg_1634[17]), .Y(n11383) );
  OAI21X1 U14529 ( .A(n5995), .B(n10036), .C(n10011), .Y(n11386) );
  AOI21X1 U14530 ( .A(n10037), .B(n10010), .C(
        CircularBuffer_len_write_assig_reg_1634[18]), .Y(n11385) );
  AOI21X1 U14531 ( .A(n11386), .B(CircularBuffer_head_i_read_ass_reg_1624[18]), 
        .C(n5336), .Y(n11388) );
  AOI21X1 U14532 ( .A(n10038), .B(n5996), .C(
        CircularBuffer_len_write_assig_reg_1634[19]), .Y(n11387) );
  OAI21X1 U14533 ( .A(n5996), .B(n10038), .C(n10009), .Y(n11390) );
  AOI21X1 U14534 ( .A(n10039), .B(n10008), .C(
        CircularBuffer_len_write_assig_reg_1634[20]), .Y(n11389) );
  AOI21X1 U14535 ( .A(n11390), .B(CircularBuffer_head_i_read_ass_reg_1624[20]), 
        .C(n5337), .Y(n11392) );
  AOI21X1 U14536 ( .A(n10040), .B(n5997), .C(
        CircularBuffer_len_write_assig_reg_1634[21]), .Y(n11391) );
  OAI21X1 U14537 ( .A(n5997), .B(n10040), .C(n10007), .Y(n11394) );
  AOI21X1 U14538 ( .A(n10041), .B(n10006), .C(
        CircularBuffer_len_write_assig_reg_1634[22]), .Y(n11393) );
  AOI21X1 U14539 ( .A(n11394), .B(CircularBuffer_head_i_read_ass_reg_1624[22]), 
        .C(n5338), .Y(n11396) );
  AOI21X1 U14540 ( .A(n10042), .B(n5998), .C(
        CircularBuffer_len_write_assig_reg_1634[23]), .Y(n11395) );
  OAI21X1 U14541 ( .A(n5998), .B(n10042), .C(n10005), .Y(n11398) );
  AOI21X1 U14542 ( .A(n10043), .B(n10004), .C(
        CircularBuffer_len_write_assig_reg_1634[24]), .Y(n11397) );
  AOI21X1 U14543 ( .A(n11398), .B(CircularBuffer_head_i_read_ass_reg_1624[24]), 
        .C(n5339), .Y(n11400) );
  AOI21X1 U14544 ( .A(n10044), .B(n5999), .C(
        CircularBuffer_len_write_assig_reg_1634[25]), .Y(n11399) );
  OAI21X1 U14545 ( .A(n5999), .B(n10044), .C(n10003), .Y(n11402) );
  AOI21X1 U14546 ( .A(n10045), .B(n10002), .C(
        CircularBuffer_len_write_assig_reg_1634[26]), .Y(n11401) );
  AOI21X1 U14547 ( .A(n11402), .B(CircularBuffer_head_i_read_ass_reg_1624[26]), 
        .C(n5340), .Y(n11404) );
  AOI21X1 U14548 ( .A(n10046), .B(n6000), .C(
        CircularBuffer_len_write_assig_reg_1634[27]), .Y(n11403) );
  OAI21X1 U14549 ( .A(n6000), .B(n10046), .C(n10001), .Y(n11406) );
  AOI21X1 U14550 ( .A(n10047), .B(n10000), .C(
        CircularBuffer_len_write_assig_reg_1634[28]), .Y(n11405) );
  AOI21X1 U14551 ( .A(n11406), .B(CircularBuffer_head_i_read_ass_reg_1624[28]), 
        .C(n5341), .Y(n11407) );
  AOI21X1 U14552 ( .A(n10048), .B(n7850), .C(
        CircularBuffer_len_write_assig_reg_1634[29]), .Y(n11408) );
  AOI21X1 U14553 ( .A(n9999), .B(CircularBuffer_head_i_read_ass_reg_1624[29]), 
        .C(n7849), .Y(n11410) );
  AOI21X1 U14554 ( .A(n10049), .B(n7848), .C(
        CircularBuffer_len_write_assig_reg_1634[30]), .Y(n11409) );
  OAI21X1 U14555 ( .A(n7848), .B(n10049), .C(n9998), .Y(\sub_1269/carry[31] )
         );
  OAI21X1 U14556 ( .A(CircularBuffer_head_i_read_ass_1_reg_1719[5]), .B(n10578), .C(\sub_1275/carry[5] ), .Y(n11411) );
  AOI21X1 U14557 ( .A(n10578), .B(CircularBuffer_head_i_read_ass_1_reg_1719[5]), .C(n10331), .Y(n11413) );
  AOI21X1 U14558 ( .A(n10333), .B(n8095), .C(
        CircularBuffer_len_read_assign_3_reg_1711[6]), .Y(n11412) );
  OAI21X1 U14559 ( .A(n8095), .B(n10333), .C(n10330), .Y(n11414) );
  OAI21X1 U14560 ( .A(CircularBuffer_len_read_assign_3_reg_1711[7]), .B(n8243), 
        .C(n8244), .Y(n11418) );
  AOI21X1 U14561 ( .A(n10334), .B(n10329), .C(
        CircularBuffer_len_read_assign_3_reg_1711[8]), .Y(n11417) );
  AOI21X1 U14562 ( .A(n11418), .B(CircularBuffer_head_i_read_ass_1_reg_1719[8]), .C(n5342), .Y(n11420) );
  AOI21X1 U14563 ( .A(n10335), .B(n7637), .C(
        CircularBuffer_len_read_assign_3_reg_1711[9]), .Y(n11419) );
  OAI21X1 U14564 ( .A(n7637), .B(n10335), .C(n10328), .Y(n11422) );
  AOI21X1 U14565 ( .A(n10336), .B(n10327), .C(
        CircularBuffer_len_read_assign_3_reg_1711[10]), .Y(n11421) );
  AOI21X1 U14566 ( .A(n11422), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[10]), .C(n5343), .Y(n11424)
         );
  AOI21X1 U14567 ( .A(n10337), .B(n6001), .C(
        CircularBuffer_len_read_assign_3_reg_1711[11]), .Y(n11423) );
  OAI21X1 U14568 ( .A(n6001), .B(n10337), .C(n10326), .Y(n11426) );
  AOI21X1 U14569 ( .A(n10338), .B(n10325), .C(
        CircularBuffer_len_read_assign_3_reg_1711[12]), .Y(n11425) );
  AOI21X1 U14570 ( .A(n11426), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[12]), .C(n5344), .Y(n11428)
         );
  AOI21X1 U14571 ( .A(n10339), .B(n6002), .C(
        CircularBuffer_len_read_assign_3_reg_1711[13]), .Y(n11427) );
  OAI21X1 U14572 ( .A(n6002), .B(n10339), .C(n10324), .Y(n11430) );
  AOI21X1 U14573 ( .A(n10340), .B(n10323), .C(
        CircularBuffer_len_read_assign_3_reg_1711[14]), .Y(n11429) );
  AOI21X1 U14574 ( .A(n11430), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[14]), .C(n5345), .Y(n11432)
         );
  AOI21X1 U14575 ( .A(n10341), .B(n6003), .C(
        CircularBuffer_len_read_assign_3_reg_1711[15]), .Y(n11431) );
  OAI21X1 U14576 ( .A(n6003), .B(n10341), .C(n10322), .Y(n11434) );
  AOI21X1 U14577 ( .A(n10342), .B(n10321), .C(
        CircularBuffer_len_read_assign_3_reg_1711[16]), .Y(n11433) );
  AOI21X1 U14578 ( .A(n11434), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[16]), .C(n5346), .Y(n11436)
         );
  AOI21X1 U14579 ( .A(n10343), .B(n6004), .C(
        CircularBuffer_len_read_assign_3_reg_1711[17]), .Y(n11435) );
  OAI21X1 U14580 ( .A(n6004), .B(n10343), .C(n10320), .Y(n11438) );
  AOI21X1 U14581 ( .A(n10344), .B(n10319), .C(
        CircularBuffer_len_read_assign_3_reg_1711[18]), .Y(n11437) );
  AOI21X1 U14582 ( .A(n11438), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[18]), .C(n5347), .Y(n11440)
         );
  AOI21X1 U14583 ( .A(n10345), .B(n6005), .C(
        CircularBuffer_len_read_assign_3_reg_1711[19]), .Y(n11439) );
  OAI21X1 U14584 ( .A(n6005), .B(n10345), .C(n10318), .Y(n11442) );
  AOI21X1 U14585 ( .A(n10346), .B(n10317), .C(
        CircularBuffer_len_read_assign_3_reg_1711[20]), .Y(n11441) );
  AOI21X1 U14586 ( .A(n11442), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[20]), .C(n5348), .Y(n11444)
         );
  AOI21X1 U14587 ( .A(n10347), .B(n6006), .C(
        CircularBuffer_len_read_assign_3_reg_1711[21]), .Y(n11443) );
  OAI21X1 U14588 ( .A(n6006), .B(n10347), .C(n10316), .Y(n11446) );
  AOI21X1 U14589 ( .A(n10348), .B(n10315), .C(
        CircularBuffer_len_read_assign_3_reg_1711[22]), .Y(n11445) );
  AOI21X1 U14590 ( .A(n11446), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[22]), .C(n5349), .Y(n11448)
         );
  AOI21X1 U14591 ( .A(n10349), .B(n6007), .C(
        CircularBuffer_len_read_assign_3_reg_1711[23]), .Y(n11447) );
  OAI21X1 U14592 ( .A(n6007), .B(n10349), .C(n10314), .Y(n11450) );
  AOI21X1 U14593 ( .A(n10350), .B(n10313), .C(
        CircularBuffer_len_read_assign_3_reg_1711[24]), .Y(n11449) );
  AOI21X1 U14594 ( .A(n11450), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[24]), .C(n5350), .Y(n11452)
         );
  AOI21X1 U14595 ( .A(n10351), .B(n6008), .C(
        CircularBuffer_len_read_assign_3_reg_1711[25]), .Y(n11451) );
  OAI21X1 U14596 ( .A(n6008), .B(n10351), .C(n10312), .Y(n11454) );
  AOI21X1 U14597 ( .A(n10352), .B(n10311), .C(
        CircularBuffer_len_read_assign_3_reg_1711[26]), .Y(n11453) );
  AOI21X1 U14598 ( .A(n11454), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[26]), .C(n5351), .Y(n11456)
         );
  AOI21X1 U14599 ( .A(n10353), .B(n8094), .C(
        CircularBuffer_len_read_assign_3_reg_1711[27]), .Y(n11455) );
  OAI21X1 U14600 ( .A(n8094), .B(n10353), .C(n10310), .Y(n11458) );
  AOI21X1 U14601 ( .A(n10354), .B(n10309), .C(
        CircularBuffer_len_read_assign_3_reg_1711[28]), .Y(n11457) );
  AOI21X1 U14602 ( .A(n11458), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[28]), .C(n5352), .Y(n11459)
         );
  AOI21X1 U14603 ( .A(n10355), .B(n8368), .C(
        CircularBuffer_len_read_assign_3_reg_1711[29]), .Y(n11460) );
  AOI21X1 U14604 ( .A(n10308), .B(
        CircularBuffer_head_i_read_ass_1_reg_1719[29]), .C(n8367), .Y(n11462)
         );
  AOI21X1 U14605 ( .A(n10356), .B(n8366), .C(
        CircularBuffer_len_read_assign_3_reg_1711[30]), .Y(n11461) );
  OAI21X1 U14606 ( .A(n8366), .B(n10356), .C(n10307), .Y(\sub_1275/carry[31] )
         );
  XOR2X1 U14607 ( .A(\add_1319/carry[31] ), .B(recentdatapoints_len[31]), .Y(
        recentdatapoints_len_load_op_fu_556_p2[31]) );
  OAI21X1 U14608 ( .A(sum_phi_fu_311_p4[14]), .B(n9703), .C(n8326), .Y(n11463)
         );
  NAND3X1 U14609 ( .A(n11474), .B(n11464), .C(n9701), .Y(n11482) );
  OAI21X1 U14610 ( .A(sum_phi_fu_311_p4[10]), .B(n9687), .C(n8327), .Y(n11465)
         );
  NAND3X1 U14611 ( .A(n8327), .B(n9687), .C(sum_phi_fu_311_p4[10]), .Y(n11467)
         );
  OAI21X1 U14612 ( .A(VCaptureThresh_loc_reg_298[12]), .B(n10065), .C(n4830), 
        .Y(n11471) );
  NOR3X1 U14613 ( .A(n8362), .B(VCaptureThresh_loc_reg_298[9]), .C(n10064), 
        .Y(n11468) );
  NAND3X1 U14614 ( .A(n9676), .B(n5572), .C(n9686), .Y(n11470) );
  OAI21X1 U14615 ( .A(n9685), .B(n11471), .C(n4831), .Y(n11480) );
  NAND3X1 U14616 ( .A(n8326), .B(n9703), .C(sum_phi_fu_311_p4[14]), .Y(n11473)
         );
  OAI21X1 U14617 ( .A(VCaptureThresh_loc_reg_298[16]), .B(n10066), .C(n4832), 
        .Y(n11478) );
  NAND3X1 U14618 ( .A(n11474), .B(n9693), .C(sum_phi_fu_311_p4[12]), .Y(n11476) );
  NAND3X1 U14619 ( .A(n5455), .B(n5573), .C(n9702), .Y(n11477) );
  OAI21X1 U14620 ( .A(n9701), .B(n11478), .C(n4833), .Y(n11479) );
  OAI21X1 U14621 ( .A(n8063), .B(n11480), .C(n11479), .Y(n11481) );
  AOI21X1 U14622 ( .A(VCaptureThresh_loc_reg_298[9]), .B(n10064), .C(n8362), 
        .Y(n11484) );
  NAND3X1 U14623 ( .A(n9685), .B(n9692), .C(n5862), .Y(n11503) );
  AOI21X1 U14624 ( .A(VCaptureThresh_loc_reg_298[2]), .B(n10061), .C(
        VCaptureThresh_loc_reg_298[1]), .Y(n11485) );
  AOI22X1 U14625 ( .A(sum_phi_fu_311_p4[1]), .B(n9654), .C(n5740), .D(
        sum_phi_fu_311_p4[0]), .Y(n11488) );
  NAND3X1 U14626 ( .A(n8353), .B(n9657), .C(sum_phi_fu_311_p4[2]), .Y(n11486)
         );
  OAI21X1 U14627 ( .A(VCaptureThresh_loc_reg_298[4]), .B(n10062), .C(n4834), 
        .Y(n11487) );
  OAI21X1 U14628 ( .A(sum_phi_fu_311_p4[6]), .B(n9668), .C(n8339), .Y(n11498)
         );
  AOI21X1 U14629 ( .A(n5511), .B(n9656), .C(n11498), .Y(n11501) );
  OAI21X1 U14630 ( .A(sum_phi_fu_311_p4[2]), .B(n9657), .C(n8353), .Y(n11491)
         );
  OAI21X1 U14631 ( .A(sum_phi_fu_311_p4[4]), .B(n9661), .C(n11495), .Y(n11490)
         );
  AOI21X1 U14632 ( .A(n9656), .B(n11491), .C(n11490), .Y(n11500) );
  NAND3X1 U14633 ( .A(n8339), .B(n9668), .C(sum_phi_fu_311_p4[6]), .Y(n11493)
         );
  OAI21X1 U14634 ( .A(VCaptureThresh_loc_reg_298[8]), .B(n10063), .C(n4835), 
        .Y(n11494) );
  AOI22X1 U14635 ( .A(sum_phi_fu_311_p4[5]), .B(n9665), .C(n11496), .D(
        sum_phi_fu_311_p4[4]), .Y(n11497) );
  AOI22X1 U14636 ( .A(n9667), .B(n11498), .C(n5722), .D(n9667), .Y(n11499) );
  AOI21X1 U14637 ( .A(n5523), .B(n5502), .C(n5296), .Y(n11502) );
  AOI22X1 U14638 ( .A(n9675), .B(n5552), .C(n5741), .D(n9675), .Y(n11504) );
  NAND3X1 U14639 ( .A(n11532), .B(n11505), .C(n5760), .Y(n11551) );
  OAI21X1 U14640 ( .A(sum_phi_fu_311_p4[18]), .B(n9717), .C(n8338), .Y(n11535)
         );
  OAI21X1 U14641 ( .A(sum_phi_fu_311_p4[22]), .B(n9734), .C(n8346), .Y(n11542)
         );
  NAND3X1 U14642 ( .A(n11539), .B(n11506), .C(n9732), .Y(n11507) );
  OAI21X1 U14643 ( .A(sum_phi_fu_311_p4[26]), .B(n9751), .C(n8322), .Y(n11511)
         );
  OAI21X1 U14644 ( .A(sum_phi_fu_311_p4[30]), .B(n9765), .C(n7832), .Y(n11508)
         );
  NAND3X1 U14645 ( .A(n11521), .B(n11509), .C(n9763), .Y(n11528) );
  OAI21X1 U14646 ( .A(n9741), .B(sum_phi_fu_311_p4[24]), .C(n11514), .Y(n11510) );
  NOR3X1 U14647 ( .A(n11511), .B(n8376), .C(n11510), .Y(n11548) );
  NAND3X1 U14648 ( .A(n9715), .B(n9723), .C(n11548), .Y(n11550) );
  NAND3X1 U14649 ( .A(n8322), .B(n9751), .C(sum_phi_fu_311_p4[26]), .Y(n11513)
         );
  OAI21X1 U14650 ( .A(VCaptureThresh_loc_reg_298[28]), .B(n10069), .C(n4836), 
        .Y(n11518) );
  NAND3X1 U14651 ( .A(n11514), .B(n9741), .C(sum_phi_fu_311_p4[24]), .Y(n11516) );
  NAND3X1 U14652 ( .A(n5456), .B(n5574), .C(n9750), .Y(n11517) );
  OAI21X1 U14653 ( .A(n9749), .B(n11518), .C(n4837), .Y(n11527) );
  MUX2X1 U14654 ( .B(n11520), .A(n10070), .S(VCaptureThresh_loc_reg_298[31]), 
        .Y(n11522) );
  NAND3X1 U14655 ( .A(n11521), .B(n9755), .C(sum_phi_fu_311_p4[28]), .Y(n11524) );
  NAND3X1 U14656 ( .A(n5457), .B(n5575), .C(n11522), .Y(n11525) );
  OAI21X1 U14657 ( .A(n9763), .B(n9764), .C(n4838), .Y(n11526) );
  OAI21X1 U14658 ( .A(n8376), .B(n11527), .C(n11526), .Y(n11547) );
  NAND3X1 U14659 ( .A(n8338), .B(n9717), .C(sum_phi_fu_311_p4[18]), .Y(n11530)
         );
  OAI21X1 U14660 ( .A(VCaptureThresh_loc_reg_298[20]), .B(n10067), .C(n4839), 
        .Y(n11531) );
  AOI22X1 U14661 ( .A(sum_phi_fu_311_p4[17]), .B(n9713), .C(n11533), .D(
        sum_phi_fu_311_p4[16]), .Y(n11534) );
  AOI22X1 U14662 ( .A(n9716), .B(n11535), .C(n5723), .D(n9716), .Y(n11544) );
  NAND3X1 U14663 ( .A(n8346), .B(n9734), .C(sum_phi_fu_311_p4[22]), .Y(n11537)
         );
  OAI21X1 U14664 ( .A(VCaptureThresh_loc_reg_298[24]), .B(n10068), .C(n4840), 
        .Y(n11538) );
  AOI22X1 U14665 ( .A(sum_phi_fu_311_p4[21]), .B(n9730), .C(n11540), .D(
        sum_phi_fu_311_p4[20]), .Y(n11541) );
  AOI22X1 U14666 ( .A(n9733), .B(n11542), .C(n5724), .D(n9733), .Y(n11543) );
  AOI21X1 U14667 ( .A(n5512), .B(n9723), .C(n5297), .Y(n11545) );
  OAI21X1 U14668 ( .A(n11548), .B(n11547), .C(n4928), .Y(n11549) );
  OAI21X1 U14669 ( .A(n5534), .B(n5701), .C(n11549), .Y(N495) );
  OAI21X1 U14670 ( .A(p_1_cast_fu_1031_p1_31), .B(n9782), .C(n7780), .Y(n11553) );
  AOI21X1 U14671 ( .A(a_thresh[23]), .B(n9490), .C(n11553), .Y(n11557) );
  OAI21X1 U14672 ( .A(p_1_cast_fu_1031_p1_31), .B(n9779), .C(n7570), .Y(n11555) );
  AOI21X1 U14673 ( .A(a_thresh[16]), .B(n9490), .C(n11555), .Y(n11556) );
  AOI21X1 U14674 ( .A(n9490), .B(a_thresh[30]), .C(n8088), .Y(n11620) );
  OAI21X1 U14675 ( .A(p_1_cast_fu_1031_p1_31), .B(n9787), .C(n7210), .Y(n11561) );
  AOI21X1 U14676 ( .A(a_thresh[24]), .B(n9490), .C(n11561), .Y(n11562) );
  OAI21X1 U14677 ( .A(p_1_cast_fu_1031_p1[6]), .B(n9770), .C(n8315), .Y(n11564) );
  AOI21X1 U14678 ( .A(a_thresh[1]), .B(n9480), .C(a_thresh[0]), .Y(n11565) );
  AOI22X1 U14679 ( .A(p_1_cast_fu_1031_p1[1]), .B(n9766), .C(n5742), .D(
        p_1_cast_fu_1031_p1[0]), .Y(n11568) );
  NAND3X1 U14680 ( .A(n8314), .B(n9767), .C(p_1_cast_fu_1031_p1[2]), .Y(n11566) );
  OAI21X1 U14681 ( .A(a_thresh[3]), .B(n9482), .C(n4841), .Y(n11567) );
  OAI21X1 U14682 ( .A(p_1_cast_fu_1031_p1[2]), .B(n9767), .C(n8314), .Y(n11571) );
  OAI21X1 U14683 ( .A(p_1_cast_fu_1031_p1[4]), .B(n9768), .C(n11576), .Y(
        n11570) );
  AOI21X1 U14684 ( .A(n9481), .B(n11571), .C(n11570), .Y(n11572) );
  NAND3X1 U14685 ( .A(n9483), .B(n5576), .C(n5863), .Y(n11601) );
  NAND3X1 U14686 ( .A(n8315), .B(n9770), .C(p_1_cast_fu_1031_p1[6]), .Y(n11575) );
  OAI21X1 U14687 ( .A(a_thresh[7]), .B(n9485), .C(n4842), .Y(n11580) );
  NAND3X1 U14688 ( .A(n11576), .B(n9768), .C(p_1_cast_fu_1031_p1[4]), .Y(
        n11578) );
  NAND3X1 U14689 ( .A(n5459), .B(n5577), .C(n9484), .Y(n11579) );
  OAI21X1 U14690 ( .A(n9483), .B(n11580), .C(n4843), .Y(n11600) );
  OAI21X1 U14691 ( .A(p_1_cast_fu_1031_p1[14]), .B(n9775), .C(n8070), .Y(
        n11581) );
  NAND3X1 U14692 ( .A(n11592), .B(n11582), .C(n9477), .Y(n11602) );
  OAI21X1 U14693 ( .A(p_1_cast_fu_1031_p1[10]), .B(n9772), .C(n8313), .Y(
        n11583) );
  NAND3X1 U14694 ( .A(n8313), .B(n9772), .C(p_1_cast_fu_1031_p1[10]), .Y(
        n11585) );
  OAI21X1 U14695 ( .A(a_thresh[11]), .B(n9475), .C(n4844), .Y(n11589) );
  NOR3X1 U14696 ( .A(n8357), .B(a_thresh[8]), .C(n9487), .Y(n11586) );
  NAND3X1 U14697 ( .A(n9486), .B(n5578), .C(n9474), .Y(n11588) );
  OAI21X1 U14698 ( .A(n9473), .B(n11589), .C(n4845), .Y(n11598) );
  NAND3X1 U14699 ( .A(n8070), .B(n9775), .C(p_1_cast_fu_1031_p1[14]), .Y(
        n11591) );
  OAI21X1 U14700 ( .A(a_thresh[15]), .B(n9479), .C(n4846), .Y(n11596) );
  NAND3X1 U14701 ( .A(n11592), .B(n9773), .C(p_1_cast_fu_1031_p1[12]), .Y(
        n11594) );
  NAND3X1 U14702 ( .A(n5460), .B(n5579), .C(n9478), .Y(n11595) );
  OAI21X1 U14703 ( .A(n9477), .B(n11596), .C(n4847), .Y(n11597) );
  OAI21X1 U14704 ( .A(n7629), .B(n11598), .C(n11597), .Y(n11599) );
  NAND3X1 U14705 ( .A(n5458), .B(n11600), .C(n9472), .Y(n11609) );
  AOI21X1 U14706 ( .A(a_thresh[8]), .B(n9487), .C(n8357), .Y(n11604) );
  NAND3X1 U14707 ( .A(n9473), .B(n9476), .C(n5864), .Y(n11607) );
  OAI21X1 U14708 ( .A(p_1_cast_fu_1031_p1_31), .B(n9781), .C(n7056), .Y(n11606) );
  AOI21X1 U14709 ( .A(n9472), .B(n5503), .C(n11606), .Y(n11608) );
  NAND3X1 U14710 ( .A(n4690), .B(n5567), .C(n5865), .Y(n11630) );
  AOI22X1 U14711 ( .A(p_1_cast_fu_1031_p1_31), .B(n9777), .C(
        p_1_cast_fu_1031_p1_31), .D(n9776), .Y(n11612) );
  AOI22X1 U14712 ( .A(p_1_cast_fu_1031_p1_31), .B(n9778), .C(
        p_1_cast_fu_1031_p1_31), .D(n9781), .Y(n11610) );
  NAND3X1 U14713 ( .A(n5353), .B(n5580), .C(n5761), .Y(n11628) );
  AOI22X1 U14714 ( .A(p_1_cast_fu_1031_p1_31), .B(n9787), .C(
        p_1_cast_fu_1031_p1_31), .D(n9786), .Y(n11614) );
  AOI22X1 U14715 ( .A(p_1_cast_fu_1031_p1_31), .B(n9785), .C(
        p_1_cast_fu_1031_p1_31), .D(n9784), .Y(n11613) );
  MUX2X1 U14716 ( .B(a_thresh[31]), .A(n7782), .S(p_1_cast_fu_1031_p1_31), .Y(
        n11617) );
  AOI22X1 U14717 ( .A(p_1_cast_fu_1031_p1_31), .B(n9789), .C(
        p_1_cast_fu_1031_p1_31), .D(n9788), .Y(n11618) );
  OAI21X1 U14718 ( .A(n8372), .B(n9489), .C(n7585), .Y(n11621) );
  OAI21X1 U14719 ( .A(n11622), .B(n5956), .C(n11621), .Y(n11623) );
  AOI22X1 U14720 ( .A(p_1_cast_fu_1031_p1_31), .B(n9780), .C(
        p_1_cast_fu_1031_p1_31), .D(n9783), .Y(n11624) );
  NAND3X1 U14721 ( .A(n9488), .B(n5581), .C(n5762), .Y(n11627) );
  OAI21X1 U14722 ( .A(n5535), .B(n5703), .C(n4929), .Y(n11629) );
  OAI21X1 U14723 ( .A(n5549), .B(n5702), .C(n11629), .Y(N496) );
  OAI21X1 U14724 ( .A(n2273), .B(n9592), .C(n7844), .Y(n11632) );
  NAND3X1 U14725 ( .A(n11643), .B(n11633), .C(n9588), .Y(n11651) );
  OAI21X1 U14726 ( .A(n2281), .B(n9579), .C(n8078), .Y(n11634) );
  NAND3X1 U14727 ( .A(n8078), .B(n9579), .C(n2281), .Y(n11636) );
  OAI21X1 U14728 ( .A(ACaptureThresh_loc_reg_288[11]), .B(n8399), .C(n4848), 
        .Y(n11640) );
  NOR3X1 U14729 ( .A(n7633), .B(ACaptureThresh_loc_reg_288[8]), .C(n8407), .Y(
        n11637) );
  NAND3X1 U14730 ( .A(n9569), .B(n7403), .C(n9576), .Y(n11639) );
  OAI21X1 U14731 ( .A(n9575), .B(n11640), .C(n7402), .Y(n11649) );
  NAND3X1 U14732 ( .A(n7844), .B(n9592), .C(n2273), .Y(n11642) );
  OAI21X1 U14733 ( .A(ACaptureThresh_loc_reg_288[15]), .B(n8114), .C(n4849), 
        .Y(n11647) );
  NAND3X1 U14734 ( .A(n11643), .B(n9584), .C(n2277), .Y(n11645) );
  NAND3X1 U14735 ( .A(n5461), .B(n5582), .C(n9589), .Y(n11646) );
  OAI21X1 U14736 ( .A(n9588), .B(n11647), .C(n4850), .Y(n11648) );
  OAI21X1 U14737 ( .A(n5952), .B(n11649), .C(n11648), .Y(n11650) );
  AOI21X1 U14738 ( .A(ACaptureThresh_loc_reg_288[8]), .B(n8407), .C(n7633), 
        .Y(n11653) );
  NAND3X1 U14739 ( .A(n9575), .B(n5951), .C(n5866), .Y(n11672) );
  AOI21X1 U14740 ( .A(ACaptureThresh_loc_reg_288[1]), .B(n10539), .C(
        ACaptureThresh_loc_reg_288[0]), .Y(n11654) );
  AOI22X1 U14741 ( .A(CircularBuffer_len_read_assign_3_fu_1091_p3[1]), .B(
        n9550), .C(n5743), .D(n2301), .Y(n11657) );
  NAND3X1 U14742 ( .A(n8352), .B(n9554), .C(
        CircularBuffer_len_read_assign_3_fu_1091_p3[2]), .Y(n11655) );
  OAI21X1 U14743 ( .A(ACaptureThresh_loc_reg_288[3]), .B(n10537), .C(n4851), 
        .Y(n11656) );
  OAI21X1 U14744 ( .A(n2289), .B(n9564), .C(n7846), .Y(n11667) );
  AOI21X1 U14745 ( .A(n5513), .B(n9552), .C(n11667), .Y(n11670) );
  OAI21X1 U14746 ( .A(CircularBuffer_len_read_assign_3_fu_1091_p3[2]), .B(
        n9554), .C(n8352), .Y(n11660) );
  OAI21X1 U14747 ( .A(CircularBuffer_len_read_assign_3_fu_1091_p3[4]), .B(
        n9558), .C(n11664), .Y(n11659) );
  AOI21X1 U14748 ( .A(n9552), .B(n11660), .C(n11659), .Y(n11669) );
  NAND3X1 U14749 ( .A(n7846), .B(n9564), .C(n2289), .Y(n11662) );
  OAI21X1 U14750 ( .A(ACaptureThresh_loc_reg_288[7]), .B(n8112), .C(n4852), 
        .Y(n11663) );
  AOI22X1 U14751 ( .A(n2291), .B(n9560), .C(n11665), .D(
        CircularBuffer_len_read_assign_3_fu_1091_p3[4]), .Y(n11666) );
  AOI22X1 U14752 ( .A(n9562), .B(n11667), .C(n5725), .D(n9562), .Y(n11668) );
  AOI21X1 U14753 ( .A(n5524), .B(n5504), .C(n5298), .Y(n11671) );
  AOI22X1 U14754 ( .A(n9568), .B(n5553), .C(n5744), .D(n9568), .Y(n11673) );
  NAND3X1 U14755 ( .A(n11701), .B(n11674), .C(n5763), .Y(n11720) );
  OAI21X1 U14756 ( .A(n2265), .B(n9604), .C(n5967), .Y(n11704) );
  OAI21X1 U14757 ( .A(n2257), .B(n9618), .C(n8086), .Y(n11711) );
  NAND3X1 U14758 ( .A(n11708), .B(n11675), .C(n9614), .Y(n11676) );
  OAI21X1 U14759 ( .A(n2249), .B(n9632), .C(n5968), .Y(n11680) );
  OAI21X1 U14760 ( .A(n2238), .B(n9644), .C(n8324), .Y(n11677) );
  NAND3X1 U14761 ( .A(n11690), .B(n11678), .C(n9640), .Y(n11697) );
  OAI21X1 U14762 ( .A(n9624), .B(n2253), .C(n11683), .Y(n11679) );
  NOR3X1 U14763 ( .A(n11680), .B(n6010), .C(n11679), .Y(n11717) );
  NAND3X1 U14764 ( .A(n9600), .B(n9608), .C(n11717), .Y(n11719) );
  NAND3X1 U14765 ( .A(n5968), .B(n9632), .C(n2249), .Y(n11682) );
  OAI21X1 U14766 ( .A(ACaptureThresh_loc_reg_288[27]), .B(n7646), .C(n4853), 
        .Y(n11687) );
  NAND3X1 U14767 ( .A(n11683), .B(n9624), .C(n2253), .Y(n11685) );
  NAND3X1 U14768 ( .A(n5462), .B(n5583), .C(n9629), .Y(n11686) );
  OAI21X1 U14769 ( .A(n9628), .B(n11687), .C(n4854), .Y(n11696) );
  NAND3X1 U14770 ( .A(n8324), .B(n9644), .C(n2238), .Y(n11689) );
  OAI21X1 U14771 ( .A(n2401), .B(n9646), .C(n4855), .Y(n11694) );
  NAND3X1 U14772 ( .A(n11690), .B(n9636), .C(n2245), .Y(n11692) );
  NAND3X1 U14773 ( .A(n5463), .B(n5584), .C(n9641), .Y(n11693) );
  OAI21X1 U14774 ( .A(n9640), .B(n11694), .C(n4856), .Y(n11695) );
  OAI21X1 U14775 ( .A(n6010), .B(n11696), .C(n11695), .Y(n11716) );
  NAND3X1 U14776 ( .A(n5967), .B(n9604), .C(n2265), .Y(n11699) );
  OAI21X1 U14777 ( .A(ACaptureThresh_loc_reg_288[19]), .B(n7864), .C(n4857), 
        .Y(n11700) );
  AOI22X1 U14778 ( .A(n2267), .B(n9598), .C(n11702), .D(n2269), .Y(n11703) );
  AOI22X1 U14779 ( .A(n9601), .B(n11704), .C(n5726), .D(n9601), .Y(n11713) );
  NAND3X1 U14780 ( .A(n8086), .B(n9618), .C(n2257), .Y(n11706) );
  OAI21X1 U14781 ( .A(ACaptureThresh_loc_reg_288[23]), .B(n8401), .C(n4858), 
        .Y(n11707) );
  AOI22X1 U14782 ( .A(n2259), .B(n9612), .C(n11709), .D(n2261), .Y(n11710) );
  AOI22X1 U14783 ( .A(n9615), .B(n11711), .C(n5727), .D(n9615), .Y(n11712) );
  AOI21X1 U14784 ( .A(n5514), .B(n9608), .C(n5299), .Y(n11714) );
  OAI21X1 U14785 ( .A(n11717), .B(n11716), .C(n4930), .Y(n11718) );
  OAI21X1 U14786 ( .A(n5536), .B(n5704), .C(n11718), .Y(N497) );
  OAI21X1 U14787 ( .A(sum_1_phi_fu_379_p4[14]), .B(n9594), .C(n8332), .Y(
        n11721) );
  NAND3X1 U14788 ( .A(n11732), .B(n11722), .C(n9354), .Y(n11740) );
  OAI21X1 U14789 ( .A(sum_1_phi_fu_379_p4[10]), .B(n9581), .C(n8333), .Y(
        n11723) );
  NAND3X1 U14790 ( .A(n8333), .B(n9581), .C(sum_1_phi_fu_379_p4[10]), .Y(
        n11725) );
  OAI21X1 U14791 ( .A(ACaptureThresh_loc_reg_288[12]), .B(n9363), .C(n4859), 
        .Y(n11729) );
  NOR3X1 U14792 ( .A(n8361), .B(ACaptureThresh_loc_reg_288[9]), .C(n9368), .Y(
        n11726) );
  NAND3X1 U14793 ( .A(n9366), .B(n5585), .C(n9362), .Y(n11728) );
  OAI21X1 U14794 ( .A(n9361), .B(n11729), .C(n4860), .Y(n11738) );
  NAND3X1 U14795 ( .A(n8332), .B(n9594), .C(sum_1_phi_fu_379_p4[14]), .Y(
        n11731) );
  OAI21X1 U14796 ( .A(ACaptureThresh_loc_reg_288[16]), .B(n9356), .C(n4861), 
        .Y(n11736) );
  NAND3X1 U14797 ( .A(n11732), .B(n9586), .C(sum_1_phi_fu_379_p4[12]), .Y(
        n11734) );
  NAND3X1 U14798 ( .A(n5464), .B(n5586), .C(n9355), .Y(n11735) );
  OAI21X1 U14799 ( .A(n9354), .B(n11736), .C(n4862), .Y(n11737) );
  OAI21X1 U14800 ( .A(n8067), .B(n11738), .C(n11737), .Y(n11739) );
  AOI21X1 U14801 ( .A(ACaptureThresh_loc_reg_288[9]), .B(n9368), .C(n8361), 
        .Y(n11742) );
  NAND3X1 U14802 ( .A(n9361), .B(n9353), .C(n5867), .Y(n11761) );
  AOI21X1 U14803 ( .A(ACaptureThresh_loc_reg_288[2]), .B(n9380), .C(
        ACaptureThresh_loc_reg_288[1]), .Y(n11743) );
  AOI22X1 U14804 ( .A(sum_1_phi_fu_379_p4[1]), .B(n9554), .C(n5745), .D(
        sum_1_phi_fu_379_p4[0]), .Y(n11746) );
  NAND3X1 U14805 ( .A(n8349), .B(n9556), .C(sum_1_phi_fu_379_p4[2]), .Y(n11744) );
  OAI21X1 U14806 ( .A(ACaptureThresh_loc_reg_288[4]), .B(n9377), .C(n4863), 
        .Y(n11745) );
  OAI21X1 U14807 ( .A(sum_1_phi_fu_379_p4[6]), .B(n9566), .C(n8350), .Y(n11756) );
  AOI21X1 U14808 ( .A(n5515), .B(n9376), .C(n11756), .Y(n11759) );
  OAI21X1 U14809 ( .A(sum_1_phi_fu_379_p4[2]), .B(n9556), .C(n8349), .Y(n11749) );
  OAI21X1 U14810 ( .A(sum_1_phi_fu_379_p4[4]), .B(n9560), .C(n11753), .Y(
        n11748) );
  AOI21X1 U14811 ( .A(n9376), .B(n11749), .C(n11748), .Y(n11758) );
  NAND3X1 U14812 ( .A(n8350), .B(n9566), .C(sum_1_phi_fu_379_p4[6]), .Y(n11751) );
  OAI21X1 U14813 ( .A(ACaptureThresh_loc_reg_288[8]), .B(n9371), .C(n4864), 
        .Y(n11752) );
  AOI22X1 U14814 ( .A(sum_1_phi_fu_379_p4[5]), .B(n9564), .C(n11754), .D(
        sum_1_phi_fu_379_p4[4]), .Y(n11755) );
  AOI22X1 U14815 ( .A(n9370), .B(n11756), .C(n5728), .D(n9370), .Y(n11757) );
  AOI21X1 U14816 ( .A(n5525), .B(n5505), .C(n5300), .Y(n11760) );
  AOI22X1 U14817 ( .A(n9352), .B(n5554), .C(n5746), .D(n9352), .Y(n11762) );
  NAND3X1 U14818 ( .A(n11790), .B(n11763), .C(n5764), .Y(n11809) );
  OAI21X1 U14819 ( .A(sum_1_phi_fu_379_p4[18]), .B(n9606), .C(n8343), .Y(
        n11793) );
  OAI21X1 U14820 ( .A(sum_1_phi_fu_379_p4[22]), .B(n9620), .C(n8342), .Y(
        n11800) );
  NAND3X1 U14821 ( .A(n11797), .B(n11764), .C(n9338), .Y(n11765) );
  OAI21X1 U14822 ( .A(sum_1_phi_fu_379_p4[26]), .B(n9634), .C(n8331), .Y(
        n11769) );
  OAI21X1 U14823 ( .A(sum_1_phi_fu_379_p4[30]), .B(n9646), .C(n7833), .Y(
        n11766) );
  NAND3X1 U14824 ( .A(n11779), .B(n11767), .C(n9323), .Y(n11786) );
  OAI21X1 U14825 ( .A(n9626), .B(sum_1_phi_fu_379_p4[24]), .C(n11772), .Y(
        n11768) );
  NOR3X1 U14826 ( .A(n11769), .B(n8377), .C(n11768), .Y(n11806) );
  NAND3X1 U14827 ( .A(n9345), .B(n9337), .C(n11806), .Y(n11808) );
  NAND3X1 U14828 ( .A(n8331), .B(n9634), .C(sum_1_phi_fu_379_p4[26]), .Y(
        n11771) );
  OAI21X1 U14829 ( .A(ACaptureThresh_loc_reg_288[28]), .B(n9332), .C(n4865), 
        .Y(n11776) );
  NAND3X1 U14830 ( .A(n11772), .B(n9626), .C(sum_1_phi_fu_379_p4[24]), .Y(
        n11774) );
  NAND3X1 U14831 ( .A(n5465), .B(n5587), .C(n9331), .Y(n11775) );
  OAI21X1 U14832 ( .A(n9330), .B(n11776), .C(n4866), .Y(n11785) );
  MUX2X1 U14833 ( .B(n11778), .A(n9325), .S(ACaptureThresh_loc_reg_288[31]), 
        .Y(n11780) );
  NAND3X1 U14834 ( .A(n11779), .B(n9638), .C(sum_1_phi_fu_379_p4[28]), .Y(
        n11782) );
  NAND3X1 U14835 ( .A(n5466), .B(n5588), .C(n11780), .Y(n11783) );
  OAI21X1 U14836 ( .A(n9323), .B(n9324), .C(n4867), .Y(n11784) );
  OAI21X1 U14837 ( .A(n8377), .B(n11785), .C(n11784), .Y(n11805) );
  NAND3X1 U14838 ( .A(n8343), .B(n9606), .C(sum_1_phi_fu_379_p4[18]), .Y(
        n11788) );
  OAI21X1 U14839 ( .A(ACaptureThresh_loc_reg_288[20]), .B(n9347), .C(n4868), 
        .Y(n11789) );
  AOI22X1 U14840 ( .A(sum_1_phi_fu_379_p4[17]), .B(n9604), .C(n11791), .D(
        sum_1_phi_fu_379_p4[16]), .Y(n11792) );
  AOI22X1 U14841 ( .A(n9346), .B(n11793), .C(n5729), .D(n9346), .Y(n11802) );
  NAND3X1 U14842 ( .A(n8342), .B(n9620), .C(sum_1_phi_fu_379_p4[22]), .Y(
        n11795) );
  OAI21X1 U14843 ( .A(ACaptureThresh_loc_reg_288[24]), .B(n9340), .C(n4869), 
        .Y(n11796) );
  AOI22X1 U14844 ( .A(sum_1_phi_fu_379_p4[21]), .B(n9618), .C(n11798), .D(
        sum_1_phi_fu_379_p4[20]), .Y(n11799) );
  AOI22X1 U14845 ( .A(n9339), .B(n11800), .C(n5730), .D(n9339), .Y(n11801) );
  AOI21X1 U14846 ( .A(n5516), .B(n9337), .C(n5301), .Y(n11803) );
  OAI21X1 U14847 ( .A(n11806), .B(n11805), .C(n4931), .Y(n11807) );
  OAI21X1 U14848 ( .A(n5537), .B(n5705), .C(n11807), .Y(N498) );
  OAI21X1 U14849 ( .A(VbeatDelay_new_1_reg_326[14]), .B(n10405), .C(n8329), 
        .Y(n11810) );
  NAND3X1 U14850 ( .A(n11821), .B(n11811), .C(n10403), .Y(n11829) );
  OAI21X1 U14851 ( .A(VbeatDelay_new_1_reg_326[10]), .B(n10394), .C(n8330), 
        .Y(n11812) );
  NAND3X1 U14852 ( .A(n8330), .B(n10394), .C(VbeatDelay_new_1_reg_326[10]), 
        .Y(n11814) );
  OAI21X1 U14853 ( .A(VbeatFallDelay_new_1_reg_342[11]), .B(n10480), .C(n7552), 
        .Y(n11818) );
  NOR3X1 U14854 ( .A(n8360), .B(VbeatFallDelay_new_1_reg_342[8]), .C(n10472), 
        .Y(n11815) );
  NAND3X1 U14855 ( .A(n10387), .B(n7788), .C(n10393), .Y(n11817) );
  OAI21X1 U14856 ( .A(n10392), .B(n11818), .C(n7787), .Y(n11827) );
  NAND3X1 U14857 ( .A(n8329), .B(n10405), .C(VbeatDelay_new_1_reg_326[14]), 
        .Y(n11820) );
  OAI21X1 U14858 ( .A(VbeatFallDelay_new_1_reg_342[15]), .B(n10491), .C(n4870), 
        .Y(n11825) );
  NAND3X1 U14859 ( .A(n11821), .B(n10399), .C(VbeatDelay_new_1_reg_326[12]), 
        .Y(n11823) );
  NAND3X1 U14860 ( .A(n5467), .B(n8239), .C(n10404), .Y(n11824) );
  OAI21X1 U14861 ( .A(n10403), .B(n11825), .C(n4871), .Y(n11826) );
  OAI21X1 U14862 ( .A(n8066), .B(n11827), .C(n11826), .Y(n11828) );
  AOI21X1 U14863 ( .A(VbeatFallDelay_new_1_reg_342[8]), .B(n10472), .C(n8360), 
        .Y(n11831) );
  NAND3X1 U14864 ( .A(n10392), .B(n10398), .C(n5868), .Y(n11850) );
  AOI21X1 U14865 ( .A(VbeatFallDelay_new_1_reg_342[1]), .B(n10454), .C(
        VbeatFallDelay_new_1_reg_342[0]), .Y(n11832) );
  AOI22X1 U14866 ( .A(VbeatDelay_new_1_reg_326[1]), .B(n10370), .C(n8249), .D(
        VbeatDelay_new_1_reg_326[0]), .Y(n11835) );
  NAND3X1 U14867 ( .A(n8347), .B(n10373), .C(VbeatDelay_new_1_reg_326[2]), .Y(
        n11833) );
  OAI21X1 U14868 ( .A(VbeatFallDelay_new_1_reg_342[3]), .B(n10459), .C(n4872), 
        .Y(n11834) );
  OAI21X1 U14869 ( .A(VbeatDelay_new_1_reg_326[6]), .B(n10382), .C(n8348), .Y(
        n11845) );
  AOI21X1 U14870 ( .A(n8248), .B(n10372), .C(n11845), .Y(n11848) );
  OAI21X1 U14871 ( .A(VbeatDelay_new_1_reg_326[2]), .B(n10373), .C(n8347), .Y(
        n11838) );
  OAI21X1 U14872 ( .A(VbeatDelay_new_1_reg_326[4]), .B(n10377), .C(n11842), 
        .Y(n11837) );
  AOI21X1 U14873 ( .A(n10372), .B(n11838), .C(n11837), .Y(n11847) );
  NAND3X1 U14874 ( .A(n8348), .B(n10382), .C(VbeatDelay_new_1_reg_326[6]), .Y(
        n11840) );
  OAI21X1 U14875 ( .A(VbeatFallDelay_new_1_reg_342[7]), .B(n10468), .C(n4873), 
        .Y(n11841) );
  AOI22X1 U14876 ( .A(VbeatDelay_new_1_reg_326[5]), .B(n10379), .C(n11843), 
        .D(VbeatDelay_new_1_reg_326[4]), .Y(n11844) );
  AOI22X1 U14877 ( .A(n10381), .B(n11845), .C(n7792), .D(n10381), .Y(n11846)
         );
  AOI21X1 U14878 ( .A(n5526), .B(n5506), .C(n5302), .Y(n11849) );
  AOI22X1 U14879 ( .A(n10386), .B(n5555), .C(n5747), .D(n10386), .Y(n11851) );
  NAND3X1 U14880 ( .A(n11879), .B(n11852), .C(n5765), .Y(n11898) );
  OAI21X1 U14881 ( .A(VbeatDelay_new_1_reg_326[18]), .B(n10415), .C(n8341), 
        .Y(n11882) );
  OAI21X1 U14882 ( .A(VbeatDelay_new_1_reg_326[22]), .B(n10426), .C(n8340), 
        .Y(n11889) );
  NAND3X1 U14883 ( .A(n11886), .B(n11853), .C(n10424), .Y(n11854) );
  OAI21X1 U14884 ( .A(VbeatDelay_new_1_reg_326[26]), .B(n10437), .C(n8328), 
        .Y(n11858) );
  OAI21X1 U14885 ( .A(VbeatDelay_new_1_reg_326[30]), .B(n10447), .C(n8076), 
        .Y(n11855) );
  NAND3X1 U14886 ( .A(n11868), .B(n11856), .C(n10445), .Y(n11875) );
  OAI21X1 U14887 ( .A(n10431), .B(VbeatDelay_new_1_reg_326[24]), .C(n11861), 
        .Y(n11857) );
  NOR3X1 U14888 ( .A(n11858), .B(n8375), .C(n11857), .Y(n11895) );
  NAND3X1 U14889 ( .A(n10413), .B(n10419), .C(n11895), .Y(n11897) );
  NAND3X1 U14890 ( .A(n8328), .B(n10437), .C(VbeatDelay_new_1_reg_326[26]), 
        .Y(n11860) );
  OAI21X1 U14891 ( .A(VbeatFallDelay_new_1_reg_342[27]), .B(n10523), .C(n4874), 
        .Y(n11865) );
  NAND3X1 U14892 ( .A(n11861), .B(n10431), .C(VbeatDelay_new_1_reg_326[24]), 
        .Y(n11863) );
  NAND3X1 U14893 ( .A(n5468), .B(n5589), .C(n10436), .Y(n11864) );
  OAI21X1 U14894 ( .A(n10435), .B(n11865), .C(n4875), .Y(n11874) );
  NAND3X1 U14895 ( .A(n8076), .B(n10447), .C(VbeatDelay_new_1_reg_326[30]), 
        .Y(n11867) );
  OAI21X1 U14896 ( .A(VbeatDelay_new_1_reg_326[31]), .B(n10449), .C(n4876), 
        .Y(n11872) );
  NAND3X1 U14897 ( .A(n11868), .B(n10441), .C(VbeatDelay_new_1_reg_326[28]), 
        .Y(n11870) );
  NAND3X1 U14898 ( .A(n5469), .B(n8003), .C(n10446), .Y(n11871) );
  OAI21X1 U14899 ( .A(n10445), .B(n11872), .C(n4877), .Y(n11873) );
  OAI21X1 U14900 ( .A(n8375), .B(n11874), .C(n11873), .Y(n11894) );
  NAND3X1 U14901 ( .A(n8341), .B(n10415), .C(VbeatDelay_new_1_reg_326[18]), 
        .Y(n11877) );
  OAI21X1 U14902 ( .A(VbeatFallDelay_new_1_reg_342[19]), .B(n10501), .C(n4878), 
        .Y(n11878) );
  AOI22X1 U14903 ( .A(VbeatDelay_new_1_reg_326[17]), .B(n10411), .C(n11880), 
        .D(VbeatDelay_new_1_reg_326[16]), .Y(n11881) );
  AOI22X1 U14904 ( .A(n10414), .B(n11882), .C(n7794), .D(n10414), .Y(n11891)
         );
  NAND3X1 U14905 ( .A(n8340), .B(n10426), .C(VbeatDelay_new_1_reg_326[22]), 
        .Y(n11884) );
  OAI21X1 U14906 ( .A(VbeatFallDelay_new_1_reg_342[23]), .B(n10512), .C(n4879), 
        .Y(n11885) );
  AOI22X1 U14907 ( .A(VbeatDelay_new_1_reg_326[21]), .B(n10422), .C(n11887), 
        .D(VbeatDelay_new_1_reg_326[20]), .Y(n11888) );
  AOI22X1 U14908 ( .A(n10425), .B(n11889), .C(n7598), .D(n10425), .Y(n11890)
         );
  AOI21X1 U14909 ( .A(n7793), .B(n10419), .C(n7597), .Y(n11892) );
  OAI21X1 U14910 ( .A(n11895), .B(n11894), .C(n4932), .Y(n11896) );
  OAI21X1 U14911 ( .A(n5538), .B(n5706), .C(n11896), .Y(N499) );
  NOR3X1 U14912 ( .A(n11899), .B(VbeatFallDelay_new_1_reg_342[24]), .C(
        VbeatFallDelay_new_1_reg_342[23]), .Y(n11902) );
  NOR3X1 U14913 ( .A(n11900), .B(VbeatFallDelay_new_1_reg_342[28]), .C(
        VbeatFallDelay_new_1_reg_342[27]), .Y(n11901) );
  NOR3X1 U14914 ( .A(VbeatFallDelay_new_1_reg_342[16]), .B(
        VbeatFallDelay_new_1_reg_342[18]), .C(VbeatFallDelay_new_1_reg_342[17]), .Y(n11903) );
  NAND3X1 U14915 ( .A(n7998), .B(n8236), .C(n11903), .Y(n11906) );
  OAI21X1 U14916 ( .A(n7790), .B(n7791), .C(n10449), .Y(n11917) );
  NOR3X1 U14917 ( .A(VbeatFallDelay_new_1_reg_342[15]), .B(
        VbeatFallDelay_new_1_reg_342[9]), .C(VbeatFallDelay_new_1_reg_342[8]), 
        .Y(n11913) );
  AOI21X1 U14918 ( .A(VbeatFallDelay_new_1_reg_342[1]), .B(
        VbeatFallDelay_new_1_reg_342[0]), .C(VbeatFallDelay_new_1_reg_342[2]), 
        .Y(n11908) );
  NAND3X1 U14919 ( .A(VbeatFallDelay_new_1_reg_342[3]), .B(n10367), .C(
        VbeatFallDelay_new_1_reg_342[4]), .Y(n11910) );
  NAND3X1 U14920 ( .A(VbeatFallDelay_new_1_reg_342[6]), .B(
        VbeatFallDelay_new_1_reg_342[5]), .C(VbeatFallDelay_new_1_reg_342[7]), 
        .Y(n11909) );
  OAI21X1 U14921 ( .A(n8005), .B(n8004), .C(n10394), .Y(n11911) );
  NOR3X1 U14922 ( .A(n11911), .B(VbeatFallDelay_new_1_reg_342[12]), .C(
        VbeatFallDelay_new_1_reg_342[11]), .Y(n11912) );
  NAND3X1 U14923 ( .A(n7589), .B(n11913), .C(n11912), .Y(n11915) );
  OAI21X1 U14924 ( .A(tmp_6_reg_1538[14]), .B(n9592), .C(n8317), .Y(n11918) );
  NAND3X1 U14925 ( .A(n11929), .B(n11919), .C(n9590), .Y(n11937) );
  OAI21X1 U14926 ( .A(tmp_6_reg_1538[10]), .B(n9579), .C(n8318), .Y(n11920) );
  NAND3X1 U14927 ( .A(n8318), .B(n9579), .C(tmp_6_reg_1538[10]), .Y(n11922) );
  OAI21X1 U14928 ( .A(ACaptureThresh_loc_reg_288[11]), .B(n10754), .C(n4880), 
        .Y(n11926) );
  NOR3X1 U14929 ( .A(n8358), .B(ACaptureThresh_loc_reg_288[8]), .C(n10751), 
        .Y(n11923) );
  NAND3X1 U14930 ( .A(n9571), .B(n7784), .C(n9578), .Y(n11925) );
  OAI21X1 U14931 ( .A(n9577), .B(n11926), .C(n7783), .Y(n11935) );
  NAND3X1 U14932 ( .A(n8317), .B(n9592), .C(tmp_6_reg_1538[14]), .Y(n11928) );
  OAI21X1 U14933 ( .A(ACaptureThresh_loc_reg_288[15]), .B(n10758), .C(n4881), 
        .Y(n11933) );
  NAND3X1 U14934 ( .A(n11929), .B(n9584), .C(tmp_6_reg_1538[12]), .Y(n11931)
         );
  NAND3X1 U14935 ( .A(n5470), .B(n8237), .C(n9591), .Y(n11932) );
  OAI21X1 U14936 ( .A(n9590), .B(n11933), .C(n4882), .Y(n11934) );
  OAI21X1 U14937 ( .A(n8064), .B(n11935), .C(n11934), .Y(n11936) );
  AOI21X1 U14938 ( .A(ACaptureThresh_loc_reg_288[8]), .B(n10751), .C(n8358), 
        .Y(n11939) );
  NAND3X1 U14939 ( .A(n9577), .B(n9583), .C(n5869), .Y(n11958) );
  AOI21X1 U14940 ( .A(ACaptureThresh_loc_reg_288[1]), .B(n10744), .C(
        ACaptureThresh_loc_reg_288[0]), .Y(n11940) );
  AOI22X1 U14941 ( .A(tmp_6_reg_1538[1]), .B(n9550), .C(n5748), .D(
        tmp_6_reg_1538[0]), .Y(n11943) );
  NAND3X1 U14942 ( .A(n8081), .B(n9554), .C(tmp_6_reg_1538[2]), .Y(n11941) );
  OAI21X1 U14943 ( .A(ACaptureThresh_loc_reg_288[3]), .B(n10746), .C(n4883), 
        .Y(n11942) );
  OAI21X1 U14944 ( .A(tmp_6_reg_1538[6]), .B(n9564), .C(n8344), .Y(n11953) );
  AOI21X1 U14945 ( .A(n5517), .B(n9553), .C(n11953), .Y(n11956) );
  OAI21X1 U14946 ( .A(tmp_6_reg_1538[2]), .B(n9554), .C(n8081), .Y(n11946) );
  OAI21X1 U14947 ( .A(tmp_6_reg_1538[4]), .B(n9558), .C(n11950), .Y(n11945) );
  AOI21X1 U14948 ( .A(n9553), .B(n11946), .C(n11945), .Y(n11955) );
  NAND3X1 U14949 ( .A(n8344), .B(n9564), .C(tmp_6_reg_1538[6]), .Y(n11948) );
  OAI21X1 U14950 ( .A(ACaptureThresh_loc_reg_288[7]), .B(n10750), .C(n4884), 
        .Y(n11949) );
  AOI22X1 U14951 ( .A(tmp_6_reg_1538[5]), .B(n9560), .C(n11951), .D(
        tmp_6_reg_1538[4]), .Y(n11952) );
  AOI22X1 U14952 ( .A(n9563), .B(n11953), .C(n8245), .D(n9563), .Y(n11954) );
  AOI21X1 U14953 ( .A(n5527), .B(n5507), .C(n5303), .Y(n11957) );
  AOI22X1 U14954 ( .A(n9570), .B(n5556), .C(n5749), .D(n9570), .Y(n11959) );
  NAND3X1 U14955 ( .A(n11987), .B(n11960), .C(n5766), .Y(n12006) );
  OAI21X1 U14956 ( .A(tmp_6_reg_1538[18]), .B(n9604), .C(n8335), .Y(n11990) );
  OAI21X1 U14957 ( .A(tmp_6_reg_1538[22]), .B(n9618), .C(n8334), .Y(n11997) );
  NAND3X1 U14958 ( .A(n11994), .B(n11961), .C(n9616), .Y(n11962) );
  OAI21X1 U14959 ( .A(tmp_6_reg_1538[26]), .B(n9632), .C(n8316), .Y(n11966) );
  OAI21X1 U14960 ( .A(tmp_6_reg_1538[30]), .B(n9644), .C(n8071), .Y(n11963) );
  NAND3X1 U14961 ( .A(n11976), .B(n11964), .C(n9642), .Y(n11983) );
  OAI21X1 U14962 ( .A(n9624), .B(tmp_6_reg_1538[24]), .C(n11969), .Y(n11965)
         );
  NOR3X1 U14963 ( .A(n11966), .B(n8373), .C(n11965), .Y(n12003) );
  NAND3X1 U14964 ( .A(n9602), .B(n9609), .C(n12003), .Y(n12005) );
  NAND3X1 U14965 ( .A(n8316), .B(n9632), .C(tmp_6_reg_1538[26]), .Y(n11968) );
  OAI21X1 U14966 ( .A(ACaptureThresh_loc_reg_288[27]), .B(n10770), .C(n4885), 
        .Y(n11973) );
  NAND3X1 U14967 ( .A(n11969), .B(n9624), .C(tmp_6_reg_1538[24]), .Y(n11971)
         );
  NAND3X1 U14968 ( .A(n5471), .B(n5590), .C(n9631), .Y(n11972) );
  OAI21X1 U14969 ( .A(n9630), .B(n11973), .C(n4886), .Y(n11982) );
  NAND3X1 U14970 ( .A(n8071), .B(n9644), .C(tmp_6_reg_1538[30]), .Y(n11975) );
  OAI21X1 U14971 ( .A(tmp_6_reg_1538[31]), .B(n9646), .C(n4887), .Y(n11980) );
  NAND3X1 U14972 ( .A(n11976), .B(n9636), .C(tmp_6_reg_1538[28]), .Y(n11978)
         );
  NAND3X1 U14973 ( .A(n5472), .B(n8000), .C(n9643), .Y(n11979) );
  OAI21X1 U14974 ( .A(n9642), .B(n11980), .C(n4888), .Y(n11981) );
  OAI21X1 U14975 ( .A(n8373), .B(n11982), .C(n11981), .Y(n12002) );
  NAND3X1 U14976 ( .A(n8335), .B(n9604), .C(tmp_6_reg_1538[18]), .Y(n11985) );
  OAI21X1 U14977 ( .A(ACaptureThresh_loc_reg_288[19]), .B(n10762), .C(n4889), 
        .Y(n11986) );
  AOI22X1 U14978 ( .A(tmp_6_reg_1538[17]), .B(n9598), .C(n11988), .D(
        tmp_6_reg_1538[16]), .Y(n11989) );
  AOI22X1 U14979 ( .A(n9603), .B(n11990), .C(n5731), .D(n9603), .Y(n11999) );
  NAND3X1 U14980 ( .A(n8334), .B(n9618), .C(tmp_6_reg_1538[22]), .Y(n11992) );
  OAI21X1 U14981 ( .A(ACaptureThresh_loc_reg_288[23]), .B(n10766), .C(n4890), 
        .Y(n11993) );
  AOI22X1 U14982 ( .A(tmp_6_reg_1538[21]), .B(n9612), .C(n11995), .D(
        tmp_6_reg_1538[20]), .Y(n11996) );
  AOI22X1 U14983 ( .A(n9617), .B(n11997), .C(n5732), .D(n9617), .Y(n11998) );
  AOI21X1 U14984 ( .A(n5518), .B(n9609), .C(n5304), .Y(n12000) );
  OAI21X1 U14985 ( .A(n12003), .B(n12002), .C(n4933), .Y(n12004) );
  OAI21X1 U14986 ( .A(n5539), .B(n5707), .C(n12004), .Y(N502) );
  OAI21X1 U14987 ( .A(tmp_7_reg_1544[14]), .B(n9699), .C(n8320), .Y(n12007) );
  NAND3X1 U14988 ( .A(n12018), .B(n12008), .C(n9695), .Y(n12026) );
  OAI21X1 U14989 ( .A(tmp_7_reg_1544[10]), .B(n9683), .C(n8321), .Y(n12009) );
  NAND3X1 U14990 ( .A(n8321), .B(n9683), .C(tmp_7_reg_1544[10]), .Y(n12011) );
  OAI21X1 U14991 ( .A(VCaptureThresh_loc_reg_298[11]), .B(n10788), .C(n4891), 
        .Y(n12015) );
  NOR3X1 U14992 ( .A(n8359), .B(VCaptureThresh_loc_reg_298[8]), .C(n10785), 
        .Y(n12012) );
  NAND3X1 U14993 ( .A(n9671), .B(n7786), .C(n9680), .Y(n12014) );
  OAI21X1 U14994 ( .A(n9679), .B(n12015), .C(n7785), .Y(n12024) );
  NAND3X1 U14995 ( .A(n8320), .B(n9699), .C(tmp_7_reg_1544[14]), .Y(n12017) );
  OAI21X1 U14996 ( .A(VCaptureThresh_loc_reg_298[15]), .B(n10792), .C(n4892), 
        .Y(n12022) );
  NAND3X1 U14997 ( .A(n12018), .B(n9690), .C(tmp_7_reg_1544[12]), .Y(n12020)
         );
  NAND3X1 U14998 ( .A(n5473), .B(n8238), .C(n9696), .Y(n12021) );
  OAI21X1 U14999 ( .A(n9695), .B(n12022), .C(n4893), .Y(n12023) );
  OAI21X1 U15000 ( .A(n8065), .B(n12024), .C(n12023), .Y(n12025) );
  AOI21X1 U15001 ( .A(VCaptureThresh_loc_reg_298[8]), .B(n10785), .C(n8359), 
        .Y(n12028) );
  NAND3X1 U15002 ( .A(n9679), .B(n9689), .C(n5870), .Y(n12047) );
  AOI21X1 U15003 ( .A(VCaptureThresh_loc_reg_298[1]), .B(n10778), .C(
        VCaptureThresh_loc_reg_298[0]), .Y(n12029) );
  AOI22X1 U15004 ( .A(tmp_7_reg_1544[1]), .B(n9650), .C(n8011), .D(
        tmp_7_reg_1544[0]), .Y(n12032) );
  NAND3X1 U15005 ( .A(n8082), .B(n9654), .C(tmp_7_reg_1544[2]), .Y(n12030) );
  OAI21X1 U15006 ( .A(VCaptureThresh_loc_reg_298[3]), .B(n10780), .C(n4894), 
        .Y(n12031) );
  OAI21X1 U15007 ( .A(tmp_7_reg_1544[6]), .B(n9665), .C(n8345), .Y(n12042) );
  AOI21X1 U15008 ( .A(n8010), .B(n9652), .C(n12042), .Y(n12045) );
  OAI21X1 U15009 ( .A(tmp_7_reg_1544[2]), .B(n9654), .C(n8082), .Y(n12035) );
  OAI21X1 U15010 ( .A(tmp_7_reg_1544[4]), .B(n9659), .C(n12039), .Y(n12034) );
  AOI21X1 U15011 ( .A(n9652), .B(n12035), .C(n12034), .Y(n12044) );
  NAND3X1 U15012 ( .A(n8345), .B(n9665), .C(tmp_7_reg_1544[6]), .Y(n12037) );
  OAI21X1 U15013 ( .A(VCaptureThresh_loc_reg_298[7]), .B(n10784), .C(n4895), 
        .Y(n12038) );
  AOI22X1 U15014 ( .A(tmp_7_reg_1544[5]), .B(n9661), .C(n12040), .D(
        tmp_7_reg_1544[4]), .Y(n12041) );
  AOI22X1 U15015 ( .A(n9663), .B(n12042), .C(n8246), .D(n9663), .Y(n12043) );
  AOI21X1 U15016 ( .A(n5528), .B(n5508), .C(n5305), .Y(n12046) );
  AOI22X1 U15017 ( .A(n9670), .B(n5557), .C(n5750), .D(n9670), .Y(n12048) );
  NAND3X1 U15018 ( .A(n12076), .B(n12049), .C(n5767), .Y(n12095) );
  OAI21X1 U15019 ( .A(tmp_7_reg_1544[18]), .B(n9713), .C(n8337), .Y(n12079) );
  OAI21X1 U15020 ( .A(tmp_7_reg_1544[22]), .B(n9730), .C(n8336), .Y(n12086) );
  NAND3X1 U15021 ( .A(n12083), .B(n12050), .C(n9726), .Y(n12051) );
  OAI21X1 U15022 ( .A(tmp_7_reg_1544[26]), .B(n9747), .C(n8319), .Y(n12055) );
  OAI21X1 U15023 ( .A(tmp_7_reg_1544[30]), .B(n9761), .C(n8072), .Y(n12052) );
  NAND3X1 U15024 ( .A(n12065), .B(n12053), .C(n9757), .Y(n12072) );
  OAI21X1 U15025 ( .A(n9738), .B(tmp_7_reg_1544[24]), .C(n12058), .Y(n12054)
         );
  NOR3X1 U15026 ( .A(n12055), .B(n8374), .C(n12054), .Y(n12092) );
  NAND3X1 U15027 ( .A(n9709), .B(n9719), .C(n12092), .Y(n12094) );
  NAND3X1 U15028 ( .A(n8319), .B(n9747), .C(tmp_7_reg_1544[26]), .Y(n12057) );
  OAI21X1 U15029 ( .A(VCaptureThresh_loc_reg_298[27]), .B(n10804), .C(n4896), 
        .Y(n12062) );
  NAND3X1 U15030 ( .A(n12058), .B(n9738), .C(tmp_7_reg_1544[24]), .Y(n12060)
         );
  NAND3X1 U15031 ( .A(n5474), .B(n5591), .C(n9744), .Y(n12061) );
  OAI21X1 U15032 ( .A(n9743), .B(n12062), .C(n4897), .Y(n12071) );
  NAND3X1 U15033 ( .A(n8072), .B(n9761), .C(tmp_7_reg_1544[30]), .Y(n12064) );
  OAI21X1 U15034 ( .A(tmp_7_reg_1544[31]), .B(n9765), .C(n4898), .Y(n12069) );
  NAND3X1 U15035 ( .A(n12065), .B(n9753), .C(tmp_7_reg_1544[28]), .Y(n12067)
         );
  NAND3X1 U15036 ( .A(n5475), .B(n8001), .C(n9758), .Y(n12068) );
  OAI21X1 U15037 ( .A(n9757), .B(n12069), .C(n4899), .Y(n12070) );
  OAI21X1 U15038 ( .A(n8374), .B(n12071), .C(n12070), .Y(n12091) );
  NAND3X1 U15039 ( .A(n8337), .B(n9713), .C(tmp_7_reg_1544[18]), .Y(n12074) );
  OAI21X1 U15040 ( .A(VCaptureThresh_loc_reg_298[19]), .B(n10796), .C(n4900), 
        .Y(n12075) );
  AOI22X1 U15041 ( .A(tmp_7_reg_1544[17]), .B(n9707), .C(n12077), .D(
        tmp_7_reg_1544[16]), .Y(n12078) );
  AOI22X1 U15042 ( .A(n9710), .B(n12079), .C(n7797), .D(n9710), .Y(n12088) );
  NAND3X1 U15043 ( .A(n8336), .B(n9730), .C(tmp_7_reg_1544[22]), .Y(n12081) );
  OAI21X1 U15044 ( .A(VCaptureThresh_loc_reg_298[23]), .B(n10800), .C(n4901), 
        .Y(n12082) );
  AOI22X1 U15045 ( .A(tmp_7_reg_1544[21]), .B(n9724), .C(n12084), .D(
        tmp_7_reg_1544[20]), .Y(n12085) );
  AOI22X1 U15046 ( .A(n9727), .B(n12086), .C(n5733), .D(n9727), .Y(n12087) );
  AOI21X1 U15047 ( .A(n7796), .B(n9719), .C(n5306), .Y(n12089) );
  OAI21X1 U15048 ( .A(n12092), .B(n12091), .C(n4934), .Y(n12093) );
  OAI21X1 U15049 ( .A(n5540), .B(n5708), .C(n12093), .Y(N505) );
  XOR2X1 U15050 ( .A(\add_1407/carry[31] ), .B(AbeatDelay[31]), .Y(
        tmp_3_fu_706_p2[31]) );
  XOR2X1 U15051 ( .A(\add_1413/carry[31] ), .B(VbeatDelay[31]), .Y(
        tmp_4_fu_716_p2[31]) );
  XOR2X1 U15052 ( .A(\add_1415/carry[31] ), .B(VbeatFallDelay[31]), .Y(
        tmp_5_fu_726_p2[31]) );
  OAI21X1 U15053 ( .A(n2766), .B(n9699), .C(n7843), .Y(n12096) );
  NAND3X1 U15054 ( .A(n12107), .B(n12097), .C(n9697), .Y(n12115) );
  OAI21X1 U15055 ( .A(n2774), .B(n9683), .C(n8077), .Y(n12098) );
  NAND3X1 U15056 ( .A(n8077), .B(n9683), .C(n2774), .Y(n12100) );
  OAI21X1 U15057 ( .A(VCaptureThresh_loc_reg_298[11]), .B(n8398), .C(n7054), 
        .Y(n12104) );
  NOR3X1 U15058 ( .A(n7632), .B(VCaptureThresh_loc_reg_298[8]), .C(n8406), .Y(
        n12101) );
  NAND3X1 U15059 ( .A(n9673), .B(n7401), .C(n9682), .Y(n12103) );
  OAI21X1 U15060 ( .A(n9681), .B(n12104), .C(n7400), .Y(n12113) );
  NAND3X1 U15061 ( .A(n7843), .B(n9699), .C(n2766), .Y(n12106) );
  OAI21X1 U15062 ( .A(VCaptureThresh_loc_reg_298[15]), .B(n8113), .C(n4902), 
        .Y(n12111) );
  NAND3X1 U15063 ( .A(n12107), .B(n9690), .C(n2770), .Y(n12109) );
  NAND3X1 U15064 ( .A(n5476), .B(n5592), .C(n9698), .Y(n12110) );
  OAI21X1 U15065 ( .A(n9697), .B(n12111), .C(n4903), .Y(n12112) );
  OAI21X1 U15066 ( .A(n5954), .B(n12113), .C(n12112), .Y(n12114) );
  AOI21X1 U15067 ( .A(VCaptureThresh_loc_reg_298[8]), .B(n8406), .C(n7632), 
        .Y(n12117) );
  NAND3X1 U15068 ( .A(n9681), .B(n5953), .C(n5871), .Y(n12136) );
  AOI21X1 U15069 ( .A(VCaptureThresh_loc_reg_298[1]), .B(n10074), .C(
        VCaptureThresh_loc_reg_298[0]), .Y(n12118) );
  AOI22X1 U15070 ( .A(CircularBuffer_len_read_assign_1_fu_778_p3[1]), .B(n9650), .C(n5751), .D(n2794), .Y(n12121) );
  NAND3X1 U15071 ( .A(n8351), .B(n9654), .C(
        CircularBuffer_len_read_assign_1_fu_778_p3[2]), .Y(n12119) );
  OAI21X1 U15072 ( .A(VCaptureThresh_loc_reg_298[3]), .B(n10072), .C(n4904), 
        .Y(n12120) );
  OAI21X1 U15073 ( .A(n2782), .B(n9665), .C(n7845), .Y(n12131) );
  AOI21X1 U15074 ( .A(n5519), .B(n9653), .C(n12131), .Y(n12134) );
  OAI21X1 U15075 ( .A(CircularBuffer_len_read_assign_1_fu_778_p3[2]), .B(n9654), .C(n8351), .Y(n12124) );
  OAI21X1 U15076 ( .A(CircularBuffer_len_read_assign_1_fu_778_p3[4]), .B(n9659), .C(n12128), .Y(n12123) );
  AOI21X1 U15077 ( .A(n9653), .B(n12124), .C(n12123), .Y(n12133) );
  NAND3X1 U15078 ( .A(n7845), .B(n9665), .C(n2782), .Y(n12126) );
  OAI21X1 U15079 ( .A(VCaptureThresh_loc_reg_298[7]), .B(n8111), .C(n4905), 
        .Y(n12127) );
  AOI22X1 U15080 ( .A(n2784), .B(n9661), .C(n12129), .D(
        CircularBuffer_len_read_assign_1_fu_778_p3[4]), .Y(n12130) );
  AOI22X1 U15081 ( .A(n9664), .B(n12131), .C(n5734), .D(n9664), .Y(n12132) );
  AOI21X1 U15082 ( .A(n5529), .B(n5509), .C(n5307), .Y(n12135) );
  AOI22X1 U15083 ( .A(n9672), .B(n5558), .C(n5752), .D(n9672), .Y(n12137) );
  NAND3X1 U15084 ( .A(n12165), .B(n12138), .C(n5768), .Y(n12184) );
  OAI21X1 U15085 ( .A(n2758), .B(n9713), .C(n5969), .Y(n12168) );
  OAI21X1 U15086 ( .A(n2750), .B(n9730), .C(n8085), .Y(n12175) );
  NAND3X1 U15087 ( .A(n12172), .B(n12139), .C(n9728), .Y(n12140) );
  OAI21X1 U15088 ( .A(n2742), .B(n9747), .C(n5970), .Y(n12144) );
  OAI21X1 U15089 ( .A(n2734), .B(n9761), .C(n8323), .Y(n12141) );
  NAND3X1 U15090 ( .A(n12154), .B(n12142), .C(n9759), .Y(n12161) );
  OAI21X1 U15091 ( .A(n9738), .B(n2746), .C(n12147), .Y(n12143) );
  NOR3X1 U15092 ( .A(n12144), .B(n6011), .C(n12143), .Y(n12181) );
  NAND3X1 U15093 ( .A(n9711), .B(n9720), .C(n12181), .Y(n12183) );
  NAND3X1 U15094 ( .A(n5970), .B(n9747), .C(n2742), .Y(n12146) );
  OAI21X1 U15095 ( .A(VCaptureThresh_loc_reg_298[27]), .B(n7645), .C(n4906), 
        .Y(n12151) );
  NAND3X1 U15096 ( .A(n12147), .B(n9738), .C(n2746), .Y(n12149) );
  NAND3X1 U15097 ( .A(n5477), .B(n5593), .C(n9746), .Y(n12150) );
  OAI21X1 U15098 ( .A(n9745), .B(n12151), .C(n4907), .Y(n12160) );
  NAND3X1 U15099 ( .A(n8323), .B(n9761), .C(n2734), .Y(n12153) );
  OAI21X1 U15100 ( .A(n2862), .B(n9765), .C(n4908), .Y(n12158) );
  NAND3X1 U15101 ( .A(n12154), .B(n9753), .C(n2738), .Y(n12156) );
  NAND3X1 U15102 ( .A(n5478), .B(n5594), .C(n9760), .Y(n12157) );
  OAI21X1 U15103 ( .A(n9759), .B(n12158), .C(n4909), .Y(n12159) );
  OAI21X1 U15104 ( .A(n6011), .B(n12160), .C(n12159), .Y(n12180) );
  NAND3X1 U15105 ( .A(n5969), .B(n9713), .C(n2758), .Y(n12163) );
  OAI21X1 U15106 ( .A(VCaptureThresh_loc_reg_298[19]), .B(n7863), .C(n4910), 
        .Y(n12164) );
  AOI22X1 U15107 ( .A(n2760), .B(n9707), .C(n12166), .D(n2762), .Y(n12167) );
  AOI22X1 U15108 ( .A(n9712), .B(n12168), .C(n5735), .D(n9712), .Y(n12177) );
  NAND3X1 U15109 ( .A(n8085), .B(n9730), .C(n2750), .Y(n12170) );
  OAI21X1 U15110 ( .A(VCaptureThresh_loc_reg_298[23]), .B(n8400), .C(n4911), 
        .Y(n12171) );
  AOI22X1 U15111 ( .A(n2752), .B(n9724), .C(n12173), .D(n2754), .Y(n12174) );
  AOI22X1 U15112 ( .A(n9729), .B(n12175), .C(n5736), .D(n9729), .Y(n12176) );
  AOI21X1 U15113 ( .A(n5520), .B(n9720), .C(n5308), .Y(n12178) );
  OAI21X1 U15114 ( .A(n12181), .B(n12180), .C(n4935), .Y(n12182) );
  OAI21X1 U15115 ( .A(n5541), .B(n5709), .C(n12182), .Y(N512) );
  OAI21X1 U15116 ( .A(p_cast_fu_688_p1_31), .B(n9523), .C(n7778), .Y(n12186)
         );
  AOI21X1 U15117 ( .A(v_thresh[23]), .B(n9540), .C(n12186), .Y(n12190) );
  OAI21X1 U15118 ( .A(p_cast_fu_688_p1_31), .B(n9520), .C(n7568), .Y(n12188)
         );
  AOI21X1 U15119 ( .A(v_thresh[16]), .B(n9540), .C(n12188), .Y(n12189) );
  AOI21X1 U15120 ( .A(n9540), .B(v_thresh[30]), .C(n8087), .Y(n12253) );
  OAI21X1 U15121 ( .A(p_cast_fu_688_p1_31), .B(n9529), .C(n7209), .Y(n12194)
         );
  AOI21X1 U15122 ( .A(v_thresh[24]), .B(n9540), .C(n12194), .Y(n12195) );
  OAI21X1 U15123 ( .A(p_cast_fu_688_p1[6]), .B(n9504), .C(n8312), .Y(n12197)
         );
  AOI21X1 U15124 ( .A(v_thresh[1]), .B(n9536), .C(v_thresh[0]), .Y(n12198) );
  AOI22X1 U15125 ( .A(p_cast_fu_688_p1[1]), .B(n9497), .C(n5753), .D(
        p_cast_fu_688_p1[0]), .Y(n12201) );
  NAND3X1 U15126 ( .A(n8311), .B(n9499), .C(p_cast_fu_688_p1[2]), .Y(n12199)
         );
  OAI21X1 U15127 ( .A(v_thresh[3]), .B(n9537), .C(n4912), .Y(n12200) );
  OAI21X1 U15128 ( .A(p_cast_fu_688_p1[2]), .B(n9499), .C(n8311), .Y(n12204)
         );
  OAI21X1 U15129 ( .A(p_cast_fu_688_p1[4]), .B(n9500), .C(n12209), .Y(n12203)
         );
  AOI21X1 U15130 ( .A(n9498), .B(n12204), .C(n12203), .Y(n12205) );
  NAND3X1 U15131 ( .A(n9502), .B(n5595), .C(n5872), .Y(n12234) );
  NAND3X1 U15132 ( .A(n8312), .B(n9504), .C(p_cast_fu_688_p1[6]), .Y(n12208)
         );
  OAI21X1 U15133 ( .A(v_thresh[7]), .B(n9538), .C(n4913), .Y(n12213) );
  NAND3X1 U15134 ( .A(n12209), .B(n9500), .C(p_cast_fu_688_p1[4]), .Y(n12211)
         );
  NAND3X1 U15135 ( .A(n5480), .B(n5596), .C(n9503), .Y(n12212) );
  OAI21X1 U15136 ( .A(n9502), .B(n12213), .C(n4914), .Y(n12233) );
  OAI21X1 U15137 ( .A(p_cast_fu_688_p1[14]), .B(n9516), .C(n8309), .Y(n12214)
         );
  NAND3X1 U15138 ( .A(n12225), .B(n12215), .C(n9514), .Y(n12235) );
  OAI21X1 U15139 ( .A(p_cast_fu_688_p1[10]), .B(n9510), .C(n8310), .Y(n12216)
         );
  NAND3X1 U15140 ( .A(n8310), .B(n9510), .C(p_cast_fu_688_p1[10]), .Y(n12218)
         );
  OAI21X1 U15141 ( .A(v_thresh[11]), .B(n9534), .C(n4915), .Y(n12222) );
  NOR3X1 U15142 ( .A(n8356), .B(v_thresh[8]), .C(n9539), .Y(n12219) );
  NAND3X1 U15143 ( .A(n9506), .B(n5597), .C(n9509), .Y(n12221) );
  OAI21X1 U15144 ( .A(n9508), .B(n12222), .C(n4916), .Y(n12231) );
  NAND3X1 U15145 ( .A(n8309), .B(n9516), .C(p_cast_fu_688_p1[14]), .Y(n12224)
         );
  OAI21X1 U15146 ( .A(v_thresh[15]), .B(n9535), .C(n4917), .Y(n12229) );
  NAND3X1 U15147 ( .A(n12225), .B(n9512), .C(p_cast_fu_688_p1[12]), .Y(n12227)
         );
  NAND3X1 U15148 ( .A(n5481), .B(n5598), .C(n9515), .Y(n12228) );
  OAI21X1 U15149 ( .A(n9514), .B(n12229), .C(n4918), .Y(n12230) );
  OAI21X1 U15150 ( .A(n8068), .B(n12231), .C(n12230), .Y(n12232) );
  NAND3X1 U15151 ( .A(n5479), .B(n12233), .C(n9505), .Y(n12242) );
  AOI21X1 U15152 ( .A(v_thresh[8]), .B(n9539), .C(n8356), .Y(n12237) );
  NAND3X1 U15153 ( .A(n9508), .B(n9511), .C(n5873), .Y(n12240) );
  OAI21X1 U15154 ( .A(p_cast_fu_688_p1_31), .B(n9522), .C(n7055), .Y(n12239)
         );
  AOI21X1 U15155 ( .A(n9505), .B(n5510), .C(n12239), .Y(n12241) );
  NAND3X1 U15156 ( .A(n4691), .B(n5568), .C(n5874), .Y(n12263) );
  AOI22X1 U15157 ( .A(p_cast_fu_688_p1_31), .B(n9518), .C(p_cast_fu_688_p1_31), 
        .D(n9517), .Y(n12245) );
  AOI22X1 U15158 ( .A(p_cast_fu_688_p1_31), .B(n9519), .C(p_cast_fu_688_p1_31), 
        .D(n9522), .Y(n12243) );
  NAND3X1 U15159 ( .A(n5354), .B(n5599), .C(n5769), .Y(n12261) );
  AOI22X1 U15160 ( .A(p_cast_fu_688_p1_31), .B(n9529), .C(p_cast_fu_688_p1_31), 
        .D(n9528), .Y(n12247) );
  AOI22X1 U15161 ( .A(p_cast_fu_688_p1_31), .B(n9527), .C(p_cast_fu_688_p1_31), 
        .D(n9526), .Y(n12246) );
  MUX2X1 U15162 ( .B(v_thresh[31]), .A(n7781), .S(p_cast_fu_688_p1_31), .Y(
        n12250) );
  AOI22X1 U15163 ( .A(p_cast_fu_688_p1_31), .B(n9531), .C(p_cast_fu_688_p1_31), 
        .D(n9530), .Y(n12251) );
  OAI21X1 U15164 ( .A(n8371), .B(n9532), .C(n7583), .Y(n12254) );
  OAI21X1 U15165 ( .A(n12255), .B(n5959), .C(n12254), .Y(n12256) );
  AOI22X1 U15166 ( .A(p_cast_fu_688_p1_31), .B(n9521), .C(p_cast_fu_688_p1_31), 
        .D(n9524), .Y(n12257) );
  NAND3X1 U15167 ( .A(n9525), .B(n5600), .C(n5770), .Y(n12260) );
  OAI21X1 U15168 ( .A(n5542), .B(n5711), .C(n4936), .Y(n12262) );
  OAI21X1 U15169 ( .A(n5550), .B(n5710), .C(n12262), .Y(N513) );
  XOR2X1 U15170 ( .A(\dp_cluster_0/add_1147_aco/carry[31] ), .B(
        \dp_cluster_0/N985 ), .Y(tmp_7_fu_511_p3[31]) );
  XOR2X1 U15171 ( .A(\dp_cluster_1/add_1107_aco/carry[31] ), .B(
        \dp_cluster_1/N953 ), .Y(tmp_6_fu_497_p3[31]) );
endmodule

